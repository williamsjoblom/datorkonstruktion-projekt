library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

-- pMem interface
entity pMem is
  port(
    pAddr : in unsigned(14 downto 0);
    pData : out unsigned(15 downto 0));
end pMem;

architecture Behavioral of pMem is

-- program Memory
type p_mem_t is array (0 to 2047) of unsigned(7 downto 0);
constant p_mem_c : p_mem_t := 
(
 x"e0"
,x"00"
,x"e8"
,x"06"
,x"9d"
,x"46"
,x"e0"
,x"e0"
,x"0f"
,x"e8"
,x"08"
,x"9d"
,x"46"
,x"e0"
,x"e0"
,x"0f"
,x"e8"
,x"09"
,x"9d"
,x"46"
,x"e0"
,x"e0"
,x"00"
,x"e8"
,x"0a"
,x"9d"
,x"46"
,x"e0"
,x"e0"
,x"fe"
,x"e8"
,x"07"
,x"9d"
,x"46"
,x"e0"
,x"9d"
,x"3c"
,x"e0"
,x"08"
,x"49"
,x"81"
,x"10"
,x"20"
,x"e0"
,x"8e"
,x"e8"
,x"00"
,x"9d"
,x"46"
,x"e0"
,x"e0"
,x"00"
,x"e8"
,x"01"
,x"9d"
,x"46"
,x"e0"
,x"7d"
,x"39"
,x"e0"
,x"09"
,x"15"
,x"20"
,x"a8"
,x"01"
,x"cd"
,x"3c"
,x"e0"
,x"a0"
,x"00"
,x"9d"
,x"3c"
,x"e0"
,x"f9"
,x"13"
,x"20"
,x"9d"
,x"3c"
,x"e0"
,x"f1"
,x"13"
,x"20"
,x"a0"
,x"00"
,x"9d"
,x"6b"
,x"e0"
,x"e8"
,x"0f"
,x"9d"
,x"85"
,x"e0"
,x"e8"
,x"00"
,x"9d"
,x"8c"
,x"e0"
,x"9d"
,x"93"
,x"e0"
,x"e8"
,x"fe"
,x"9d"
,x"9a"
,x"e0"
,x"a0"
,x"00"
,x"9d"
,x"aa"
,x"e0"
,x"e0"
,x"06"
,x"e8"
,x"00"
,x"9d"
,x"77"
,x"e0"
,x"a0"
,x"00"
,x"9d"
,x"b3"
,x"e0"
,x"f1"
,x"13"
,x"20"
,x"9d"
,x"b3"
,x"e0"
,x"f9"
,x"13"
,x"20"
,x"a0"
,x"00"
,x"e0"
,x"08"
,x"9d"
,x"77"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"09"
,x"9d"
,x"77"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"0a"
,x"9d"
,x"77"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"07"
,x"9d"
,x"77"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"07"
,x"e8"
,x"f8"
,x"9d"
,x"77"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"07"
,x"e8"
,x"ff"
,x"9d"
,x"77"
,x"e0"
,x"a0"
,x"00"
,x"09"
,x"15"
,x"20"
,x"a8"
,x"01"
,x"cd"
,x"b3"
,x"e0"
,x"a0"
,x"00"
,x"08"
,x"00"
,x"81"
,x"02"
,x"20"
,x"81"
,x"03"
,x"20"
,x"a0"
,x"00"
,x"82"
,x"40"
,x"fa"
,x"41"
,x"18"
,x"00"
,x"20"
,x"00"
,x"e0"
,x"00"
,x"0f"
,x"40"
,x"00"
,x"a8"
,x"00"
,x"bd"
,x"e1"
,x"e0"
,x"9d"
,x"e3"
,x"e0"
,x"68"
,x"00"
,x"7d"
,x"d1"
,x"e0"
,x"a0"
,x"00"
,x"84"
,x"04"
,x"20"
,x"fc"
,x"06"
,x"20"
,x"9d"
,x"13"
,x"e1"
,x"a0"
,x"00"
,x"88"
,x"00"
,x"60"
,x"04"
,x"9d"
,x"fe"
,x"e0"
,x"90"
,x"00"
,x"40"
,x"0f"
,x"9d"
,x"fe"
,x"e0"
,x"a0"
,x"00"
,x"e8"
,x"f0"
,x"a8"
,x"0a"
,x"d5"
,x"0c"
,x"e1"
,x"30"
,x"30"
,x"9d"
,x"e3"
,x"e0"
,x"a0"
,x"00"
,x"30"
,x"37"
,x"9d"
,x"e3"
,x"e0"
,x"a0"
,x"00"
,x"09"
,x"02"
,x"20"
,x"a8"
,x"4f"
,x"bd"
,x"22"
,x"e1"
,x"30"
,x"01"
,x"81"
,x"02"
,x"20"
,x"a0"
,x"00"
,x"08"
,x"00"
,x"81"
,x"02"
,x"20"
,x"09"
,x"03"
,x"20"
,x"a8"
,x"3b"
,x"bd"
,x"36"
,x"e1"
,x"30"
,x"01"
,x"81"
,x"03"
,x"20"
,x"a0"
,x"00"
,x"08"
,x"00"
,x"81"
,x"03"
,x"20"
,x"a0"
,x"00"
,x"f1"
,x"02"
,x"20"
,x"f9"
,x"03"
,x"20"
,x"a0"
,x"00"
,x"43"
,x"68"
,x"20"
,x"41"
,x"20"
,x"20"
,x"20"
,x"20"
,x"43"
,x"68"
,x"20"
,x"42"
,x"20"
,x"20"
,x"20"
,x"20"
,x"43"
,x"68"
,x"20"
,x"43"
,x"00"
,x"43"
,x"20"
,x"00"
,x"43"
,x"23"
,x"00"
,x"44"
,x"20"
,x"00"
,x"44"
,x"23"
,x"00"
,x"45"
,x"20"
,x"00"
,x"46"
,x"20"
,x"00"
,x"46"
,x"23"
,x"00"
,x"47"
,x"20"
,x"00"
,x"47"
,x"23"
,x"00"
,x"41"
,x"20"
,x"00"
,x"41"
,x"23"
,x"00"
,x"42"
,x"20"
,x"00"
,x"2d"
,x"2d"
,x"20"
,x"00"
,x"65"
,x"72"
,x"72"
,x"00"
,x"08"
,x"00"
,x"82"
,x"60"
,x"82"
,x"61"
,x"e8"
,x"0f"
,x"9d"
,x"85"
,x"e0"
,x"9d"
,x"8c"
,x"e0"
,x"9d"
,x"93"
,x"e0"
,x"e0"
,x"0b"
,x"e8"
,x"e1"
,x"08"
,x"45"
,x"9d"
,x"c7"
,x"e0"
,x"9d"
,x"3a"
,x"e4"
,x"9d"
,x"52"
,x"e4"
,x"9d"
,x"6a"
,x"e4"
,x"e0"
,x"00"
,x"e8"
,x"01"
,x"9d"
,x"3d"
,x"e1"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"e8"
,x"f8"
,x"fa"
,x"6c"
,x"9d"
,x"9a"
,x"e0"
,x"a0"
,x"00"
,x"e8"
,x"ff"
,x"fa"
,x"6c"
,x"9d"
,x"9a"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"6c"
,x"40"
,x"fe"
,x"82"
,x"6c"
,x"20"
,x"00"
,x"9d"
,x"9a"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"6c"
,x"40"
,x"fd"
,x"82"
,x"6c"
,x"20"
,x"00"
,x"9d"
,x"9a"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"6c"
,x"40"
,x"fb"
,x"82"
,x"6c"
,x"20"
,x"00"
,x"9d"
,x"9a"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"6c"
,x"48"
,x"01"
,x"82"
,x"6c"
,x"20"
,x"00"
,x"9d"
,x"9a"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"6c"
,x"48"
,x"02"
,x"82"
,x"6c"
,x"20"
,x"00"
,x"9d"
,x"9a"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"6c"
,x"48"
,x"04"
,x"82"
,x"6c"
,x"20"
,x"00"
,x"9d"
,x"9a"
,x"e0"
,x"a0"
,x"00"
,x"09"
,x"08"
,x"20"
,x"40"
,x"08"
,x"a8"
,x"00"
,x"bd"
,x"2e"
,x"e2"
,x"09"
,x"08"
,x"20"
,x"40"
,x"08"
,x"a8"
,x"00"
,x"cd"
,x"21"
,x"e2"
,x"9d"
,x"b9"
,x"e2"
,x"09"
,x"08"
,x"20"
,x"40"
,x"04"
,x"a8"
,x"00"
,x"bd"
,x"45"
,x"e2"
,x"09"
,x"08"
,x"20"
,x"40"
,x"04"
,x"a8"
,x"00"
,x"cd"
,x"38"
,x"e2"
,x"9d"
,x"ce"
,x"e2"
,x"09"
,x"08"
,x"20"
,x"40"
,x"02"
,x"a8"
,x"00"
,x"bd"
,x"5c"
,x"e2"
,x"09"
,x"08"
,x"20"
,x"40"
,x"02"
,x"a8"
,x"00"
,x"cd"
,x"4f"
,x"e2"
,x"9d"
,x"e3"
,x"e2"
,x"09"
,x"08"
,x"20"
,x"40"
,x"01"
,x"a8"
,x"00"
,x"bd"
,x"73"
,x"e2"
,x"09"
,x"08"
,x"20"
,x"40"
,x"01"
,x"a8"
,x"00"
,x"cd"
,x"66"
,x"e2"
,x"9d"
,x"f8"
,x"e2"
,x"a0"
,x"00"
,x"9d"
,x"89"
,x"e2"
,x"0a"
,x"60"
,x"58"
,x"03"
,x"10"
,x"00"
,x"0a"
,x"61"
,x"30"
,x"01"
,x"20"
,x"00"
,x"9d"
,x"3d"
,x"e1"
,x"a0"
,x"00"
,x"0a"
,x"61"
,x"a8"
,x"00"
,x"d5"
,x"97"
,x"e2"
,x"08"
,x"26"
,x"82"
,x"61"
,x"7d"
,x"a0"
,x"e2"
,x"a8"
,x"27"
,x"c5"
,x"a0"
,x"e2"
,x"08"
,x"00"
,x"82"
,x"61"
,x"0a"
,x"60"
,x"a8"
,x"00"
,x"d5"
,x"ae"
,x"e2"
,x"08"
,x"02"
,x"82"
,x"60"
,x"7d"
,x"b7"
,x"e2"
,x"a8"
,x"03"
,x"c5"
,x"b7"
,x"e2"
,x"08"
,x"00"
,x"82"
,x"60"
,x"a0"
,x"00"
,x"08"
,x"f0"
,x"84"
,x"06"
,x"20"
,x"0a"
,x"61"
,x"38"
,x"01"
,x"82"
,x"61"
,x"9d"
,x"75"
,x"e2"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"08"
,x"f0"
,x"84"
,x"06"
,x"20"
,x"0a"
,x"60"
,x"30"
,x"01"
,x"82"
,x"60"
,x"9d"
,x"75"
,x"e2"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"08"
,x"f0"
,x"84"
,x"06"
,x"20"
,x"0a"
,x"61"
,x"30"
,x"01"
,x"82"
,x"61"
,x"9d"
,x"75"
,x"e2"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"9d"
,x"b1"
,x"e4"
,x"a0"
,x"00"
,x"08"
,x"f0"
,x"84"
,x"06"
,x"20"
,x"0a"
,x"60"
,x"38"
,x"01"
,x"82"
,x"60"
,x"9d"
,x"75"
,x"e2"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"9d"
,x"5d"
,x"e5"
,x"a8"
,x"01"
,x"bd"
,x"1c"
,x"e3"
,x"a0"
,x"00"
,x"9d"
,x"42"
,x"e5"
,x"a8"
,x"01"
,x"c5"
,x"1c"
,x"e3"
,x"58"
,x"04"
,x"82"
,x"6f"
,x"9d"
,x"42"
,x"e5"
,x"4a"
,x"6f"
,x"20"
,x"00"
,x"e2"
,x"61"
,x"0a"
,x"60"
,x"a8"
,x"00"
,x"bd"
,x"42"
,x"e3"
,x"a8"
,x"01"
,x"bd"
,x"4b"
,x"e3"
,x"a8"
,x"02"
,x"bd"
,x"54"
,x"e3"
,x"fb"
,x"00"
,x"10"
,x"9d"
,x"3a"
,x"e4"
,x"7d"
,x"5a"
,x"e3"
,x"fb"
,x"00"
,x"11"
,x"9d"
,x"52"
,x"e4"
,x"7d"
,x"5a"
,x"e3"
,x"fb"
,x"00"
,x"12"
,x"9d"
,x"6a"
,x"e4"
,x"9d"
,x"75"
,x"e2"
,x"a0"
,x"00"
,x"9d"
,x"17"
,x"e2"
,x"9d"
,x"12"
,x"e3"
,x"a0"
,x"00"
,x"a8"
,x"ff"
,x"bd"
,x"7e"
,x"e3"
,x"88"
,x"00"
,x"60"
,x"04"
,x"9d"
,x"fe"
,x"e0"
,x"90"
,x"00"
,x"e0"
,x"f0"
,x"40"
,x"0f"
,x"9d"
,x"89"
,x"e3"
,x"a0"
,x"00"
,x"e0"
,x"f0"
,x"e8"
,x"e1"
,x"08"
,x"7e"
,x"9d"
,x"c7"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"00"
,x"cd"
,x"97"
,x"e3"
,x"e8"
,x"e1"
,x"08"
,x"5a"
,x"9d"
,x"c7"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"01"
,x"cd"
,x"a5"
,x"e3"
,x"e8"
,x"e1"
,x"08"
,x"5d"
,x"9d"
,x"c7"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"02"
,x"cd"
,x"b3"
,x"e3"
,x"e8"
,x"e1"
,x"08"
,x"60"
,x"9d"
,x"c7"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"03"
,x"cd"
,x"c1"
,x"e3"
,x"e8"
,x"e1"
,x"08"
,x"63"
,x"9d"
,x"c7"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"04"
,x"cd"
,x"cf"
,x"e3"
,x"e8"
,x"e1"
,x"08"
,x"66"
,x"9d"
,x"c7"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"05"
,x"cd"
,x"dd"
,x"e3"
,x"e8"
,x"e1"
,x"08"
,x"69"
,x"9d"
,x"c7"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"06"
,x"cd"
,x"eb"
,x"e3"
,x"e8"
,x"e1"
,x"08"
,x"6c"
,x"9d"
,x"c7"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"07"
,x"cd"
,x"f9"
,x"e3"
,x"e8"
,x"e1"
,x"08"
,x"6f"
,x"9d"
,x"c7"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"08"
,x"cd"
,x"07"
,x"e4"
,x"e8"
,x"e1"
,x"08"
,x"72"
,x"9d"
,x"c7"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"09"
,x"cd"
,x"15"
,x"e4"
,x"e8"
,x"e1"
,x"08"
,x"75"
,x"9d"
,x"c7"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"0a"
,x"cd"
,x"23"
,x"e4"
,x"e8"
,x"e1"
,x"08"
,x"78"
,x"9d"
,x"c7"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"0b"
,x"cd"
,x"31"
,x"e4"
,x"e8"
,x"e1"
,x"08"
,x"7b"
,x"9d"
,x"c7"
,x"e0"
,x"a0"
,x"00"
,x"e8"
,x"e1"
,x"08"
,x"82"
,x"9d"
,x"c7"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"00"
,x"e8"
,x"01"
,x"9d"
,x"3d"
,x"e1"
,x"e8"
,x"10"
,x"08"
,x"00"
,x"9d"
,x"82"
,x"e4"
,x"9d"
,x"75"
,x"e2"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"e0"
,x"08"
,x"e8"
,x"01"
,x"9d"
,x"3d"
,x"e1"
,x"e8"
,x"11"
,x"08"
,x"00"
,x"9d"
,x"82"
,x"e4"
,x"9d"
,x"75"
,x"e2"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"e0"
,x"10"
,x"e8"
,x"01"
,x"9d"
,x"3d"
,x"e1"
,x"e8"
,x"12"
,x"08"
,x"00"
,x"9d"
,x"82"
,x"e4"
,x"9d"
,x"75"
,x"e2"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"82"
,x"50"
,x"fa"
,x"51"
,x"e0"
,x"00"
,x"18"
,x"00"
,x"88"
,x"00"
,x"0f"
,x"50"
,x"00"
,x"9d"
,x"67"
,x"e3"
,x"90"
,x"00"
,x"10"
,x"00"
,x"09"
,x"02"
,x"20"
,x"38"
,x"03"
,x"81"
,x"02"
,x"20"
,x"09"
,x"03"
,x"20"
,x"30"
,x"01"
,x"81"
,x"03"
,x"20"
,x"68"
,x"00"
,x"18"
,x"00"
,x"a8"
,x"27"
,x"cd"
,x"88"
,x"e4"
,x"a0"
,x"00"
,x"08"
,x"00"
,x"88"
,x"00"
,x"9d"
,x"b7"
,x"e1"
,x"90"
,x"00"
,x"10"
,x"00"
,x"88"
,x"00"
,x"9d"
,x"e9"
,x"e4"
,x"90"
,x"00"
,x"10"
,x"00"
,x"88"
,x"00"
,x"9d"
,x"00"
,x"e5"
,x"90"
,x"00"
,x"10"
,x"00"
,x"88"
,x"00"
,x"9d"
,x"17"
,x"e5"
,x"90"
,x"00"
,x"30"
,x"01"
,x"a8"
,x"27"
,x"bd"
,x"e4"
,x"e4"
,x"88"
,x"00"
,x"9d"
,x"2e"
,x"e5"
,x"7d"
,x"b5"
,x"e4"
,x"9d"
,x"c0"
,x"e1"
,x"a0"
,x"00"
,x"e3"
,x"00"
,x"10"
,x"18"
,x"00"
,x"a8"
,x"ff"
,x"cd"
,x"f8"
,x"e4"
,x"9d"
,x"f0"
,x"e1"
,x"a0"
,x"00"
,x"9d"
,x"b3"
,x"e0"
,x"f1"
,x"10"
,x"20"
,x"a0"
,x"00"
,x"e3"
,x"00"
,x"11"
,x"18"
,x"00"
,x"a8"
,x"ff"
,x"cd"
,x"0f"
,x"e5"
,x"9d"
,x"fd"
,x"e1"
,x"a0"
,x"00"
,x"9d"
,x"b3"
,x"e0"
,x"f1"
,x"11"
,x"20"
,x"a0"
,x"00"
,x"e3"
,x"00"
,x"12"
,x"18"
,x"00"
,x"a8"
,x"ff"
,x"cd"
,x"26"
,x"e5"
,x"9d"
,x"0a"
,x"e2"
,x"a0"
,x"00"
,x"9d"
,x"b3"
,x"e0"
,x"f1"
,x"12"
,x"20"
,x"a0"
,x"00"
,x"08"
,x"14"
,x"e0"
,x"fa"
,x"88"
,x"00"
,x"9d"
,x"6f"
,x"e5"
,x"90"
,x"00"
,x"38"
,x"01"
,x"a8"
,x"00"
,x"cd"
,x"32"
,x"e5"
,x"a0"
,x"00"
,x"09"
,x"09"
,x"20"
,x"40"
,x"f0"
,x"a8"
,x"00"
,x"cd"
,x"42"
,x"e5"
,x"e1"
,x"09"
,x"20"
,x"09"
,x"09"
,x"20"
,x"40"
,x"f0"
,x"a8"
,x"00"
,x"bd"
,x"4f"
,x"e5"
,x"18"
,x"00"
,x"a0"
,x"00"
,x"09"
,x"09"
,x"20"
,x"40"
,x"f0"
,x"a8"
,x"00"
,x"bd"
,x"6b"
,x"e5"
,x"08"
,x"00"
,x"a0"
,x"00"
,x"08"
,x"01"
,x"a0"
,x"00"
,x"e8"
,x"ff"
,x"28"
,x"00"
,x"38"
,x"01"
,x"20"
,x"00"
,x"a8"
,x"00"
,x"cd"
,x"71"
,x"e5"
,x"18"
,x"00"
,x"38"
,x"01"
,x"10"
,x"00"
,x"a8"
,x"00"
,x"cd"
,x"6f"
,x"e5"
,x"a0"
,x"00"
,x"77"
,x"0b"
,x"a6"
,x"47"
,x"ec"
,x"97"
,x"47"
,x"fb"
,x"b3"
,x"70"
,x"30"
,x"f4"
,x"00"
,x"00"
,x"00"
,x"00"
,x"bb"
,x"85"
,x"53"
,x"23"
,x"f6"
,x"cb"
,x"a3"
,x"7d"
,x"59"
,x"38"
,x"18"
,x"fa"
,x"00"
,x"00"
,x"00"
,x"00"
,x"dd"
,x"c2"
,x"a9"
,x"91"
,x"7b"
,x"65"
,x"51"
,x"3e"
,x"2c"
,x"1c"
,x"0c"
,x"fd"
,x"00"
,x"00"
,x"00"
,x"00"
,x"ee"
,x"e1"
,x"d4"
,x"c8"
,x"bd"
,x"b2"
,x"a8"
,x"9f"
,x"96"
,x"8e"
,x"86"
,x"7e"
,x"00"
,x"00"
,x"00"
,x"00"
,x"77"
,x"70"
,x"6a"
,x"64"
,x"5e"
,x"59"
,x"54"
,x"4f"
,x"4b"
,x"47"
,x"43"
,x"3f"
,x"00"
,x"00"
,x"00"
,x"00"
,x"3b"
,x"38"
,x"35"
,x"32"
,x"2f"
,x"2c"
,x"2a"
,x"27"
,x"25"
,x"23"
,x"21"
,x"1f"
,x"00"
,x"00"
,x"00"
,x"00"
,x"1d"
,x"1c"
,x"1a"
,x"19"
,x"17"
,x"16"
,x"15"
,x"13"
,x"12"
,x"11"
,x"10"
,x"0f"
,x"00"
,x"00"
,x"00"
,x"00"
,x"0e"
,x"0e"
,x"0d"
,x"0c"
,x"0b"
,x"0b"
,x"0a"
,x"09"
,x"09"
,x"08"
,x"08"
,x"07"
,x"00"
,x"00"
,x"00"
,x"00"
,x"07"
,x"07"
,x"06"
,x"06"
,x"05"
,x"05"
,x"05"
,x"04"
,x"04"
,x"04"
,x"04"
,x"03"
,x"00"
,x"00"
,x"00"
,x"00"
,x"07"
,x"07"
,x"06"
,x"06"
,x"05"
,x"05"
,x"05"
,x"04"
,x"04"
,x"04"
,x"04"
,x"03"
,x"00"
,x"00"
,x"00"
,x"00"
,x"03"
,x"03"
,x"03"
,x"03"
,x"02"
,x"02"
,x"02"
,x"02"
,x"02"
,x"02"
,x"02"
,x"01"
,x"00"
,x"00"
,x"00"
,x"00"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"e0"
);


  signal p_mem : p_mem_t := p_mem_c;


begin  -- pMem
  pData <= p_mem(to_integer(pAddr(10 downto 0) + 1)) & p_mem(to_integer(pAddr(10 downto 0)));

end Behavioral;

