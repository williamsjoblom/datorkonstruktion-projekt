library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

-- pMem interface
entity pMem is
  port(
    pAddr : in unsigned(14 downto 0);
    pData : out unsigned(15 downto 0));
end pMem;

architecture Behavioral of pMem is

-- program Memory
type p_mem_t is array (0 to 4095) of unsigned(7 downto 0);
constant p_mem_c : p_mem_t := 
(
 x"9d"
,x"9b"
,x"e0"
,x"9d"
,x"0f"
,x"e0"
,x"9d"
,x"8f"
,x"e3"
,x"9d"
,x"f4"
,x"e5"
,x"7d"
,x"09"
,x"e0"
,x"9d"
,x"2d"
,x"e0"
,x"9d"
,x"92"
,x"e0"
,x"e0"
,x"06"
,x"e8"
,x"00"
,x"9d"
,x"25"
,x"e0"
,x"e0"
,x"0d"
,x"e8"
,x"0c"
,x"9d"
,x"25"
,x"e0"
,x"a0"
,x"00"
,x"9d"
,x"4a"
,x"e0"
,x"9d"
,x"3a"
,x"e0"
,x"a0"
,x"00"
,x"08"
,x"00"
,x"81"
,x"01"
,x"20"
,x"9d"
,x"64"
,x"e0"
,x"9d"
,x"5a"
,x"e0"
,x"a0"
,x"00"
,x"f9"
,x"00"
,x"20"
,x"08"
,x"fe"
,x"81"
,x"01"
,x"20"
,x"9d"
,x"64"
,x"e0"
,x"9d"
,x"5a"
,x"e0"
,x"a0"
,x"00"
,x"f1"
,x"00"
,x"20"
,x"08"
,x"ff"
,x"81"
,x"01"
,x"20"
,x"9d"
,x"64"
,x"e0"
,x"9d"
,x"5a"
,x"e0"
,x"a0"
,x"00"
,x"08"
,x"04"
,x"81"
,x"01"
,x"20"
,x"9d"
,x"64"
,x"e0"
,x"a0"
,x"00"
,x"08"
,x"14"
,x"38"
,x"01"
,x"cd"
,x"66"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"08"
,x"9d"
,x"25"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"09"
,x"9d"
,x"25"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"0a"
,x"9d"
,x"25"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"07"
,x"9d"
,x"25"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"07"
,x"e8"
,x"f8"
,x"9d"
,x"25"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"07"
,x"e8"
,x"ff"
,x"9d"
,x"25"
,x"e0"
,x"a0"
,x"00"
,x"08"
,x"00"
,x"81"
,x"02"
,x"20"
,x"81"
,x"03"
,x"20"
,x"a0"
,x"00"
,x"82"
,x"40"
,x"fa"
,x"41"
,x"18"
,x"00"
,x"20"
,x"00"
,x"e0"
,x"00"
,x"0f"
,x"40"
,x"00"
,x"a8"
,x"00"
,x"bd"
,x"bf"
,x"e0"
,x"9d"
,x"c1"
,x"e0"
,x"68"
,x"00"
,x"7d"
,x"af"
,x"e0"
,x"a0"
,x"00"
,x"84"
,x"04"
,x"20"
,x"fc"
,x"06"
,x"20"
,x"9d"
,x"f1"
,x"e0"
,x"a0"
,x"00"
,x"88"
,x"00"
,x"60"
,x"04"
,x"9d"
,x"dc"
,x"e0"
,x"90"
,x"00"
,x"40"
,x"0f"
,x"9d"
,x"dc"
,x"e0"
,x"a0"
,x"00"
,x"e8"
,x"f0"
,x"a8"
,x"0a"
,x"d5"
,x"ea"
,x"e0"
,x"30"
,x"30"
,x"9d"
,x"c1"
,x"e0"
,x"a0"
,x"00"
,x"30"
,x"37"
,x"9d"
,x"c1"
,x"e0"
,x"a0"
,x"00"
,x"09"
,x"02"
,x"20"
,x"a8"
,x"4f"
,x"bd"
,x"00"
,x"e1"
,x"30"
,x"01"
,x"81"
,x"02"
,x"20"
,x"a0"
,x"00"
,x"08"
,x"00"
,x"81"
,x"02"
,x"20"
,x"09"
,x"03"
,x"20"
,x"a8"
,x"3b"
,x"bd"
,x"14"
,x"e1"
,x"30"
,x"01"
,x"81"
,x"03"
,x"20"
,x"a0"
,x"00"
,x"08"
,x"00"
,x"81"
,x"03"
,x"20"
,x"a0"
,x"00"
,x"f1"
,x"02"
,x"20"
,x"f9"
,x"03"
,x"20"
,x"a0"
,x"00"
,x"43"
,x"68"
,x"20"
,x"41"
,x"20"
,x"20"
,x"20"
,x"20"
,x"43"
,x"68"
,x"20"
,x"42"
,x"20"
,x"20"
,x"20"
,x"20"
,x"43"
,x"68"
,x"20"
,x"43"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"00"
,x"20"
,x"28"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"29"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"29"
,x"20"
,x"20"
,x"28"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"29"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"29"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"2a"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"00"
,x"20"
,x"29"
,x"5c"
,x"20"
,x"29"
,x"20"
,x"20"
,x"28"
,x"20"
,x"2f"
,x"28"
,x"20"
,x"20"
,x"20"
,x"28"
,x"20"
,x"2f"
,x"28"
,x"20"
,x"20"
,x"29"
,x"5c"
,x"20"
,x"29"
,x"20"
,x"20"
,x"20"
,x"28"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"28"
,x"20"
,x"20"
,x"20"
,x"28"
,x"20"
,x"2f"
,x"28"
,x"20"
,x"20"
,x"20"
,x"28"
,x"20"
,x"2f"
,x"28"
,x"20"
,x"20"
,x"20"
,x"28"
,x"20"
,x"20"
,x"60"
,x"20"
,x"20"
,x"20"
,x"20"
,x"00"
,x"28"
,x"28"
,x"29"
,x"2f"
,x"28"
,x"20"
,x"20"
,x"29"
,x"5c"
,x"28"
,x"29"
,x"29"
,x"20"
,x"20"
,x"29"
,x"5c"
,x"28"
,x"29"
,x"29"
,x"28"
,x"28"
,x"29"
,x"2f"
,x"28"
,x"20"
,x"20"
,x"20"
,x"29"
,x"5c"
,x"20"
,x"20"
,x"20"
,x"20"
,x"28"
,x"20"
,x"29"
,x"5c"
,x"20"
,x"20"
,x"29"
,x"5c"
,x"28"
,x"29"
,x"29"
,x"20"
,x"20"
,x"29"
,x"5c"
,x"28"
,x"29"
,x"29"
,x"20"
,x"20"
,x"29"
,x"5c"
,x"29"
,x"29"
,x"28"
,x"20"
,x"20"
,x"20"
,x"00"
,x"20"
,x"2f"
,x"28"
,x"5f"
,x"29"
,x"29"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"5c"
,x"20"
,x"20"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"5c"
,x"20"
,x"20"
,x"2f"
,x"28"
,x"5f"
,x"29"
,x"29"
,x"28"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"20"
,x"20"
,x"20"
,x"29"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"5c"
,x"20"
,x"20"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"5c"
,x"20"
,x"20"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"28"
,x"29"
,x"5c"
,x"20"
,x"20"
,x"00"
,x"28"
,x"5f"
,x"29"
,x"29"
,x"20"
,x"20"
,x"20"
,x"20"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"20"
,x"20"
,x"5f"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"28"
,x"5f"
,x"29"
,x"29"
,x"20"
,x"20"
,x"29"
,x"5c"
,x"5f"
,x"5f"
,x"5f"
,x"20"
,x"20"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"5f"
,x"20"
,x"20"
,x"20"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"20"
,x"20"
,x"20"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"20"
,x"28"
,x"5f"
,x"28"
,x"29"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"20"
,x"00"
,x"2f"
,x"20"
,x"5f"
,x"5f"
,x"7c"
,x"20"
,x"20"
,x"2f"
,x"20"
,x"5f"
,x"20"
,x"5c"
,x"20"
,x"7c"
,x"20"
,x"5c"
,x"7c"
,x"20"
,x"7c"
,x"7c"
,x"5f"
,x"20"
,x"5f"
,x"7c"
,x"28"
,x"28"
,x"2f"
,x"20"
,x"5f"
,x"5f"
,x"7c"
,x"20"
,x"20"
,x"7c"
,x"20"
,x"5f"
,x"20"
,x"29"
,x"20"
,x"2f"
,x"20"
,x"5f"
,x"20"
,x"5c"
,x"20"
,x"20"
,x"2f"
,x"20"
,x"5f"
,x"20"
,x"5c"
,x"20"
,x"7c"
,x"20"
,x"20"
,x"5c"
,x"2f"
,x"20"
,x"20"
,x"7c"
,x"20"
,x"00"
,x"5c"
,x"5f"
,x"5f"
,x"20"
,x"5c"
,x"20"
,x"7c"
,x"20"
,x"28"
,x"5f"
,x"29"
,x"20"
,x"7c"
,x"7c"
,x"20"
,x"2e"
,x"60"
,x"20"
,x"7c"
,x"20"
,x"7c"
,x"20"
,x"7c"
,x"20"
,x"20"
,x"7c"
,x"20"
,x"28"
,x"5f"
,x"5f"
,x"20"
,x"20"
,x"20"
,x"7c"
,x"20"
,x"5f"
,x"20"
,x"5c"
,x"7c"
,x"20"
,x"28"
,x"5f"
,x"29"
,x"20"
,x"7c"
,x"7c"
,x"20"
,x"28"
,x"5f"
,x"29"
,x"20"
,x"7c"
,x"7c"
,x"20"
,x"7c"
,x"5c"
,x"2f"
,x"7c"
,x"20"
,x"7c"
,x"20"
,x"00"
,x"7c"
,x"5f"
,x"5f"
,x"5f"
,x"2f"
,x"20"
,x"20"
,x"5c"
,x"5f"
,x"5f"
,x"5f"
,x"2f"
,x"20"
,x"7c"
,x"5f"
,x"7c"
,x"5c"
,x"5f"
,x"7c"
,x"7c"
,x"5f"
,x"5f"
,x"5f"
,x"7c"
,x"20"
,x"20"
,x"5c"
,x"5f"
,x"5f"
,x"5f"
,x"7c"
,x"20"
,x"20"
,x"7c"
,x"5f"
,x"5f"
,x"5f"
,x"2f"
,x"20"
,x"5c"
,x"5f"
,x"5f"
,x"5f"
,x"2f"
,x"20"
,x"20"
,x"5c"
,x"5f"
,x"5f"
,x"5f"
,x"2f"
,x"20"
,x"7c"
,x"5f"
,x"7c"
,x"20"
,x"20"
,x"7c"
,x"5f"
,x"7c"
,x"20"
,x"00"
,x"43"
,x"20"
,x"00"
,x"43"
,x"23"
,x"00"
,x"44"
,x"20"
,x"00"
,x"44"
,x"23"
,x"00"
,x"45"
,x"20"
,x"00"
,x"46"
,x"20"
,x"00"
,x"46"
,x"23"
,x"00"
,x"47"
,x"20"
,x"00"
,x"47"
,x"23"
,x"00"
,x"41"
,x"20"
,x"00"
,x"41"
,x"23"
,x"00"
,x"42"
,x"20"
,x"00"
,x"2d"
,x"2d"
,x"20"
,x"00"
,x"65"
,x"72"
,x"00"
,x"08"
,x"00"
,x"82"
,x"60"
,x"82"
,x"61"
,x"08"
,x"01"
,x"82"
,x"6d"
,x"e8"
,x"0f"
,x"9d"
,x"6d"
,x"e0"
,x"9d"
,x"74"
,x"e0"
,x"9d"
,x"7b"
,x"e0"
,x"9d"
,x"46"
,x"e7"
,x"e0"
,x"0b"
,x"e8"
,x"e1"
,x"08"
,x"23"
,x"9d"
,x"a5"
,x"e0"
,x"9d"
,x"cf"
,x"e6"
,x"9d"
,x"e7"
,x"e6"
,x"9d"
,x"ff"
,x"e6"
,x"e0"
,x"00"
,x"e8"
,x"01"
,x"9d"
,x"1b"
,x"e1"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"9d"
,x"ca"
,x"e3"
,x"a0"
,x"00"
,x"e0"
,x"09"
,x"e8"
,x"29"
,x"9d"
,x"1b"
,x"e1"
,x"e0"
,x"e0"
,x"e8"
,x"e1"
,x"08"
,x"74"
,x"9d"
,x"a5"
,x"e0"
,x"e0"
,x"09"
,x"e8"
,x"2a"
,x"9d"
,x"1b"
,x"e1"
,x"e0"
,x"e0"
,x"e8"
,x"e1"
,x"08"
,x"b2"
,x"9d"
,x"a5"
,x"e0"
,x"e0"
,x"09"
,x"e8"
,x"2b"
,x"9d"
,x"1b"
,x"e1"
,x"e0"
,x"e0"
,x"e8"
,x"e1"
,x"08"
,x"f0"
,x"9d"
,x"a5"
,x"e0"
,x"e0"
,x"09"
,x"e8"
,x"2c"
,x"9d"
,x"1b"
,x"e1"
,x"e0"
,x"e0"
,x"e8"
,x"e2"
,x"08"
,x"2e"
,x"9d"
,x"a5"
,x"e0"
,x"e0"
,x"09"
,x"e8"
,x"2d"
,x"9d"
,x"1b"
,x"e1"
,x"e0"
,x"e0"
,x"e8"
,x"e2"
,x"08"
,x"6c"
,x"9d"
,x"a5"
,x"e0"
,x"e0"
,x"09"
,x"e8"
,x"2e"
,x"9d"
,x"1b"
,x"e1"
,x"e0"
,x"f0"
,x"e8"
,x"e2"
,x"08"
,x"aa"
,x"9d"
,x"a5"
,x"e0"
,x"e0"
,x"09"
,x"e8"
,x"2f"
,x"9d"
,x"1b"
,x"e1"
,x"e0"
,x"f0"
,x"e8"
,x"e2"
,x"08"
,x"e8"
,x"9d"
,x"a5"
,x"e0"
,x"e0"
,x"09"
,x"e8"
,x"30"
,x"9d"
,x"1b"
,x"e1"
,x"e0"
,x"f0"
,x"e8"
,x"e3"
,x"08"
,x"26"
,x"9d"
,x"a5"
,x"e0"
,x"a0"
,x"00"
,x"e8"
,x"f8"
,x"fa"
,x"6c"
,x"9d"
,x"82"
,x"e0"
,x"a0"
,x"00"
,x"e8"
,x"ff"
,x"fa"
,x"6c"
,x"9d"
,x"82"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"6c"
,x"40"
,x"fe"
,x"82"
,x"6c"
,x"20"
,x"00"
,x"9d"
,x"82"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"6c"
,x"40"
,x"fd"
,x"82"
,x"6c"
,x"20"
,x"00"
,x"9d"
,x"82"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"6c"
,x"40"
,x"fb"
,x"82"
,x"6c"
,x"20"
,x"00"
,x"9d"
,x"82"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"6c"
,x"48"
,x"01"
,x"82"
,x"6c"
,x"20"
,x"00"
,x"9d"
,x"82"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"6c"
,x"48"
,x"02"
,x"82"
,x"6c"
,x"20"
,x"00"
,x"9d"
,x"82"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"6c"
,x"48"
,x"04"
,x"82"
,x"6c"
,x"20"
,x"00"
,x"9d"
,x"82"
,x"e0"
,x"a0"
,x"00"
,x"09"
,x"08"
,x"20"
,x"40"
,x"08"
,x"a8"
,x"00"
,x"bd"
,x"c3"
,x"e4"
,x"09"
,x"08"
,x"20"
,x"40"
,x"08"
,x"a8"
,x"00"
,x"cd"
,x"b6"
,x"e4"
,x"9d"
,x"4e"
,x"e5"
,x"09"
,x"08"
,x"20"
,x"40"
,x"04"
,x"a8"
,x"00"
,x"bd"
,x"da"
,x"e4"
,x"09"
,x"08"
,x"20"
,x"40"
,x"04"
,x"a8"
,x"00"
,x"cd"
,x"cd"
,x"e4"
,x"9d"
,x"63"
,x"e5"
,x"09"
,x"08"
,x"20"
,x"40"
,x"02"
,x"a8"
,x"00"
,x"bd"
,x"f1"
,x"e4"
,x"09"
,x"08"
,x"20"
,x"40"
,x"02"
,x"a8"
,x"00"
,x"cd"
,x"e4"
,x"e4"
,x"9d"
,x"78"
,x"e5"
,x"09"
,x"08"
,x"20"
,x"40"
,x"01"
,x"a8"
,x"00"
,x"bd"
,x"08"
,x"e5"
,x"09"
,x"08"
,x"20"
,x"40"
,x"01"
,x"a8"
,x"00"
,x"cd"
,x"fb"
,x"e4"
,x"9d"
,x"8d"
,x"e5"
,x"a0"
,x"00"
,x"9d"
,x"1e"
,x"e5"
,x"0a"
,x"60"
,x"58"
,x"03"
,x"10"
,x"00"
,x"0a"
,x"61"
,x"30"
,x"01"
,x"20"
,x"00"
,x"9d"
,x"1b"
,x"e1"
,x"a0"
,x"00"
,x"0a"
,x"61"
,x"a8"
,x"00"
,x"d5"
,x"2c"
,x"e5"
,x"08"
,x"26"
,x"82"
,x"61"
,x"7d"
,x"35"
,x"e5"
,x"a8"
,x"27"
,x"c5"
,x"35"
,x"e5"
,x"08"
,x"00"
,x"82"
,x"61"
,x"0a"
,x"60"
,x"a8"
,x"00"
,x"d5"
,x"43"
,x"e5"
,x"08"
,x"02"
,x"82"
,x"60"
,x"7d"
,x"4c"
,x"e5"
,x"a8"
,x"03"
,x"c5"
,x"4c"
,x"e5"
,x"08"
,x"00"
,x"82"
,x"60"
,x"a0"
,x"00"
,x"08"
,x"f0"
,x"84"
,x"06"
,x"20"
,x"0a"
,x"61"
,x"38"
,x"01"
,x"82"
,x"61"
,x"9d"
,x"0a"
,x"e5"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"08"
,x"f0"
,x"84"
,x"06"
,x"20"
,x"0a"
,x"60"
,x"30"
,x"01"
,x"82"
,x"60"
,x"9d"
,x"0a"
,x"e5"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"08"
,x"f0"
,x"84"
,x"06"
,x"20"
,x"0a"
,x"61"
,x"30"
,x"01"
,x"82"
,x"61"
,x"9d"
,x"0a"
,x"e5"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"9d"
,x"5e"
,x"e7"
,x"a0"
,x"00"
,x"08"
,x"f0"
,x"84"
,x"06"
,x"20"
,x"0a"
,x"60"
,x"38"
,x"01"
,x"82"
,x"60"
,x"9d"
,x"0a"
,x"e5"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"9d"
,x"7c"
,x"e8"
,x"a8"
,x"01"
,x"bd"
,x"b1"
,x"e5"
,x"a0"
,x"00"
,x"9d"
,x"61"
,x"e8"
,x"a8"
,x"01"
,x"c5"
,x"b1"
,x"e5"
,x"58"
,x"04"
,x"82"
,x"6f"
,x"9d"
,x"61"
,x"e8"
,x"4a"
,x"6f"
,x"20"
,x"00"
,x"e2"
,x"61"
,x"0a"
,x"60"
,x"a8"
,x"00"
,x"bd"
,x"d7"
,x"e5"
,x"a8"
,x"01"
,x"bd"
,x"e0"
,x"e5"
,x"a8"
,x"02"
,x"bd"
,x"e9"
,x"e5"
,x"fb"
,x"00"
,x"10"
,x"9d"
,x"cf"
,x"e6"
,x"7d"
,x"ef"
,x"e5"
,x"fb"
,x"00"
,x"11"
,x"9d"
,x"e7"
,x"e6"
,x"7d"
,x"ef"
,x"e5"
,x"fb"
,x"00"
,x"12"
,x"9d"
,x"ff"
,x"e6"
,x"9d"
,x"0a"
,x"e5"
,x"a0"
,x"00"
,x"9d"
,x"ac"
,x"e4"
,x"9d"
,x"a7"
,x"e5"
,x"a0"
,x"00"
,x"a8"
,x"ff"
,x"bd"
,x"13"
,x"e6"
,x"88"
,x"00"
,x"60"
,x"04"
,x"9d"
,x"dc"
,x"e0"
,x"90"
,x"00"
,x"e0"
,x"f0"
,x"40"
,x"0f"
,x"9d"
,x"1e"
,x"e6"
,x"a0"
,x"00"
,x"e0"
,x"f0"
,x"e8"
,x"e3"
,x"08"
,x"88"
,x"9d"
,x"a5"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"00"
,x"cd"
,x"2c"
,x"e6"
,x"e8"
,x"e3"
,x"08"
,x"64"
,x"9d"
,x"a5"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"01"
,x"cd"
,x"3a"
,x"e6"
,x"e8"
,x"e3"
,x"08"
,x"67"
,x"9d"
,x"a5"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"02"
,x"cd"
,x"48"
,x"e6"
,x"e8"
,x"e3"
,x"08"
,x"6a"
,x"9d"
,x"a5"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"03"
,x"cd"
,x"56"
,x"e6"
,x"e8"
,x"e3"
,x"08"
,x"6d"
,x"9d"
,x"a5"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"04"
,x"cd"
,x"64"
,x"e6"
,x"e8"
,x"e3"
,x"08"
,x"70"
,x"9d"
,x"a5"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"05"
,x"cd"
,x"72"
,x"e6"
,x"e8"
,x"e3"
,x"08"
,x"73"
,x"9d"
,x"a5"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"06"
,x"cd"
,x"80"
,x"e6"
,x"e8"
,x"e3"
,x"08"
,x"76"
,x"9d"
,x"a5"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"07"
,x"cd"
,x"8e"
,x"e6"
,x"e8"
,x"e3"
,x"08"
,x"79"
,x"9d"
,x"a5"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"08"
,x"cd"
,x"9c"
,x"e6"
,x"e8"
,x"e3"
,x"08"
,x"7c"
,x"9d"
,x"a5"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"09"
,x"cd"
,x"aa"
,x"e6"
,x"e8"
,x"e3"
,x"08"
,x"7f"
,x"9d"
,x"a5"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"0a"
,x"cd"
,x"b8"
,x"e6"
,x"e8"
,x"e3"
,x"08"
,x"82"
,x"9d"
,x"a5"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"0b"
,x"cd"
,x"c6"
,x"e6"
,x"e8"
,x"e3"
,x"08"
,x"85"
,x"9d"
,x"a5"
,x"e0"
,x"a0"
,x"00"
,x"e8"
,x"e3"
,x"08"
,x"8c"
,x"9d"
,x"a5"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"00"
,x"e8"
,x"01"
,x"9d"
,x"1b"
,x"e1"
,x"e8"
,x"10"
,x"08"
,x"00"
,x"9d"
,x"17"
,x"e7"
,x"9d"
,x"0a"
,x"e5"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"e0"
,x"08"
,x"e8"
,x"01"
,x"9d"
,x"1b"
,x"e1"
,x"e8"
,x"11"
,x"08"
,x"00"
,x"9d"
,x"17"
,x"e7"
,x"9d"
,x"0a"
,x"e5"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"e0"
,x"10"
,x"e8"
,x"01"
,x"9d"
,x"1b"
,x"e1"
,x"e8"
,x"12"
,x"08"
,x"00"
,x"9d"
,x"17"
,x"e7"
,x"9d"
,x"0a"
,x"e5"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"82"
,x"50"
,x"fa"
,x"51"
,x"e0"
,x"00"
,x"18"
,x"00"
,x"88"
,x"00"
,x"0f"
,x"50"
,x"00"
,x"9d"
,x"fc"
,x"e5"
,x"90"
,x"00"
,x"10"
,x"00"
,x"09"
,x"02"
,x"20"
,x"38"
,x"03"
,x"81"
,x"02"
,x"20"
,x"09"
,x"03"
,x"20"
,x"30"
,x"01"
,x"81"
,x"03"
,x"20"
,x"68"
,x"00"
,x"18"
,x"00"
,x"a8"
,x"27"
,x"cd"
,x"1d"
,x"e7"
,x"a0"
,x"00"
,x"e0"
,x"00"
,x"08"
,x"ff"
,x"83"
,x"00"
,x"10"
,x"83"
,x"00"
,x"11"
,x"83"
,x"00"
,x"12"
,x"68"
,x"00"
,x"18"
,x"00"
,x"a8"
,x"27"
,x"cd"
,x"48"
,x"e7"
,x"a0"
,x"00"
,x"08"
,x"00"
,x"88"
,x"00"
,x"9d"
,x"4c"
,x"e4"
,x"90"
,x"00"
,x"10"
,x"00"
,x"9d"
,x"1a"
,x"e8"
,x"88"
,x"00"
,x"9d"
,x"99"
,x"e7"
,x"90"
,x"00"
,x"10"
,x"00"
,x"88"
,x"00"
,x"9d"
,x"c4"
,x"e7"
,x"90"
,x"00"
,x"10"
,x"00"
,x"88"
,x"00"
,x"9d"
,x"ef"
,x"e7"
,x"90"
,x"00"
,x"30"
,x"01"
,x"a8"
,x"27"
,x"bd"
,x"94"
,x"e7"
,x"88"
,x"00"
,x"9d"
,x"4d"
,x"e8"
,x"7d"
,x"62"
,x"e7"
,x"9d"
,x"55"
,x"e4"
,x"a0"
,x"00"
,x"0b"
,x"00"
,x"10"
,x"38"
,x"10"
,x"10"
,x"00"
,x"a8"
,x"ff"
,x"cd"
,x"aa"
,x"e7"
,x"9d"
,x"85"
,x"e4"
,x"a0"
,x"00"
,x"0b"
,x"a8"
,x"e8"
,x"82"
,x"6a"
,x"0b"
,x"38"
,x"e9"
,x"82"
,x"6b"
,x"e0"
,x"00"
,x"ea"
,x"6a"
,x"9d"
,x"25"
,x"e0"
,x"e0"
,x"01"
,x"ea"
,x"6b"
,x"9d"
,x"25"
,x"e0"
,x"a0"
,x"00"
,x"e3"
,x"00"
,x"11"
,x"38"
,x"10"
,x"18"
,x"00"
,x"a8"
,x"ff"
,x"cd"
,x"d5"
,x"e7"
,x"9d"
,x"92"
,x"e4"
,x"a0"
,x"00"
,x"0b"
,x"a8"
,x"e8"
,x"82"
,x"6a"
,x"0b"
,x"38"
,x"e9"
,x"82"
,x"6b"
,x"e0"
,x"02"
,x"ea"
,x"6a"
,x"9d"
,x"25"
,x"e0"
,x"e0"
,x"03"
,x"ea"
,x"6b"
,x"9d"
,x"25"
,x"e0"
,x"a0"
,x"00"
,x"e3"
,x"00"
,x"12"
,x"38"
,x"10"
,x"18"
,x"00"
,x"a8"
,x"ff"
,x"cd"
,x"00"
,x"e8"
,x"9d"
,x"9f"
,x"e4"
,x"a0"
,x"00"
,x"0b"
,x"a8"
,x"e8"
,x"82"
,x"6a"
,x"0b"
,x"38"
,x"e9"
,x"82"
,x"6b"
,x"e0"
,x"04"
,x"ea"
,x"6a"
,x"9d"
,x"25"
,x"e0"
,x"e0"
,x"05"
,x"ea"
,x"6b"
,x"9d"
,x"25"
,x"e0"
,x"a0"
,x"00"
,x"18"
,x"00"
,x"88"
,x"00"
,x"9d"
,x"42"
,x"e8"
,x"e8"
,x"f0"
,x"08"
,x"20"
,x"9d"
,x"c1"
,x"e0"
,x"90"
,x"00"
,x"88"
,x"00"
,x"10"
,x"00"
,x"30"
,x"01"
,x"82"
,x"6d"
,x"9d"
,x"42"
,x"e8"
,x"e8"
,x"f0"
,x"08"
,x"3c"
,x"9d"
,x"c1"
,x"e0"
,x"90"
,x"00"
,x"10"
,x"00"
,x"a0"
,x"00"
,x"0a"
,x"6d"
,x"20"
,x"00"
,x"e0"
,x"14"
,x"9d"
,x"1b"
,x"e1"
,x"a0"
,x"00"
,x"08"
,x"0a"
,x"e0"
,x"fa"
,x"88"
,x"00"
,x"9d"
,x"8e"
,x"e8"
,x"90"
,x"00"
,x"38"
,x"01"
,x"a8"
,x"00"
,x"cd"
,x"51"
,x"e8"
,x"a0"
,x"00"
,x"09"
,x"09"
,x"20"
,x"40"
,x"f0"
,x"a8"
,x"00"
,x"cd"
,x"61"
,x"e8"
,x"e1"
,x"09"
,x"20"
,x"09"
,x"09"
,x"20"
,x"40"
,x"f0"
,x"a8"
,x"00"
,x"bd"
,x"6e"
,x"e8"
,x"18"
,x"00"
,x"a0"
,x"00"
,x"09"
,x"09"
,x"20"
,x"40"
,x"f0"
,x"a8"
,x"00"
,x"bd"
,x"8a"
,x"e8"
,x"08"
,x"00"
,x"a0"
,x"00"
,x"08"
,x"01"
,x"a0"
,x"00"
,x"e8"
,x"ff"
,x"28"
,x"00"
,x"38"
,x"01"
,x"20"
,x"00"
,x"a8"
,x"00"
,x"cd"
,x"90"
,x"e8"
,x"18"
,x"00"
,x"38"
,x"01"
,x"10"
,x"00"
,x"a8"
,x"00"
,x"cd"
,x"8e"
,x"e8"
,x"a0"
,x"00"
,x"77"
,x"0b"
,x"a6"
,x"47"
,x"ec"
,x"97"
,x"47"
,x"fb"
,x"b3"
,x"70"
,x"30"
,x"f4"
,x"00"
,x"00"
,x"00"
,x"00"
,x"bb"
,x"85"
,x"53"
,x"23"
,x"f6"
,x"cb"
,x"a3"
,x"7d"
,x"59"
,x"38"
,x"18"
,x"fa"
,x"00"
,x"00"
,x"00"
,x"00"
,x"dd"
,x"c2"
,x"a9"
,x"91"
,x"7b"
,x"65"
,x"51"
,x"3e"
,x"2c"
,x"1c"
,x"0c"
,x"fd"
,x"00"
,x"00"
,x"00"
,x"00"
,x"ee"
,x"e1"
,x"d4"
,x"c8"
,x"bd"
,x"b2"
,x"a8"
,x"9f"
,x"96"
,x"8e"
,x"86"
,x"7e"
,x"00"
,x"00"
,x"00"
,x"00"
,x"77"
,x"70"
,x"6a"
,x"64"
,x"5e"
,x"59"
,x"54"
,x"4f"
,x"4b"
,x"47"
,x"43"
,x"3f"
,x"00"
,x"00"
,x"00"
,x"00"
,x"3b"
,x"38"
,x"35"
,x"32"
,x"2f"
,x"2c"
,x"2a"
,x"27"
,x"25"
,x"23"
,x"21"
,x"1f"
,x"00"
,x"00"
,x"00"
,x"00"
,x"1d"
,x"1c"
,x"1a"
,x"19"
,x"17"
,x"16"
,x"15"
,x"13"
,x"12"
,x"11"
,x"10"
,x"0f"
,x"00"
,x"00"
,x"00"
,x"00"
,x"0e"
,x"0e"
,x"0d"
,x"0c"
,x"0b"
,x"0b"
,x"0a"
,x"09"
,x"09"
,x"08"
,x"08"
,x"07"
,x"00"
,x"00"
,x"00"
,x"00"
,x"07"
,x"07"
,x"06"
,x"06"
,x"05"
,x"05"
,x"05"
,x"04"
,x"04"
,x"04"
,x"04"
,x"03"
,x"00"
,x"00"
,x"00"
,x"00"
,x"07"
,x"07"
,x"06"
,x"06"
,x"05"
,x"05"
,x"05"
,x"04"
,x"04"
,x"04"
,x"04"
,x"03"
,x"00"
,x"00"
,x"00"
,x"00"
,x"03"
,x"03"
,x"03"
,x"03"
,x"02"
,x"02"
,x"02"
,x"02"
,x"02"
,x"02"
,x"02"
,x"01"
,x"00"
,x"00"
,x"00"
,x"00"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"e0"
);


  signal p_mem : p_mem_t := p_mem_c;


begin  -- pMem
  pData <= p_mem(to_integer(pAddr(11 downto 0) + 1)) & p_mem(to_integer(pAddr(11 downto 0)));

end Behavioral;

