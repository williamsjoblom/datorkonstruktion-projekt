library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

-- uMem interface
entity uMem is
  port (
    uAddr : in unsigned(7 downto 0);
    uData : out unsigned(28 downto 0));
end uMem;

architecture Behavioral of uMem is

-- micro Memory
type u_mem_t is array (0 to 255) of unsigned(28 downto 0);
constant u_mem_c : u_mem_t :=
  -- ALU__TB___FB__PC_LC_SEQ__uAddr
   -- Fetch
  (b"0000_0011_1111_0_00_00_0000_00000000", -- ASR := PC
   b"0000_0010_0001_1_00_00_0000_00000000", -- IR := PM, PC++
   -- E-A Calculation
   b"0000_0000_0000_0_00_00_0010_00000000", -- uPC := K2
   -- Immediate Addressing
   b"0000_0011_1110_1_00_00_0001_00000000", -- ASR := PC, PC++, uPC := K1
   -- Absolute Addressing
   b"0000_0010_1110_1_00_00_0000_00000000", -- ASR := PM, PC++
   b"0000_0000_0000_1_00_00_0001_00000000", -- PC++, uPC := K1 
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000"
   );

signal u_mem : u_mem_t := u_mem_c;

begin  -- Behavioral
  uData <= u_mem(to_integer(uAddr));

end Behavioral;
