library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

-- uMem interface
entity uMem is
  port (
    uAddr : in unsigned(7 downto 0);
    uData : out unsigned(28 downto 0));
end uMem;

architecture Behavioral of uMem is


-- micro Memory
type u_mem_t is array (0 to 255) of unsigned(28 downto 0);
constant u_mem_c : u_mem_t :=
  -- ALU__TB___FB__PC_LC_ST_SEQ__uAddr
   -- Fetch
  (b"0000_0011_1110_0_00_00_0000_00000000", -- ASR := PC
   b"0000_0010_0001_1_00_00_0000_00000000", -- IR := PM, PC++
   -- E-A Calculation
   b"0000_0000_0000_0_00_00_0010_00000000", -- uPC := K2
   -- Immediate Addressing: LDA #10
   b"0000_0011_1110_1_00_00_0001_00000000", -- ASR := PC, PC++, uPC := K1
   -- Absolute Addressing: JMP $FF77
   b"0000_0011_1110_1_00_00_0000_00000000", -- ASR := PC, PC++
   b"0000_0010_1110_1_00_00_0000_00000000", -- ASR := PM, PC++
   b"0000_0000_0000_1_00_00_0001_00000000", -- PC++, uPC := K1
   -- ZP Absolute Addressing: JMP $33
   b"0000_0011_1110_1_00_00_0000_00000000", -- ASR := PC, PC++
   b"0000_0010_1110_1_00_00_0000_00000000", -- ASR := PM, PC++
   b"0000_0000_1111_0_00_00_0001_00000000", -- ASRmsb := 0, uPC := K1
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   -- NOP
   b"0000_0000_0000_0_00_00_0011_00000000", -- uPC := 0
   -- LDA
   b"0001_0010_0000_0_00_00_0011_00000000", -- A := PM, uPC := 0
   -- TAX
   b"0000_0111_1000_0_00_00_0011_00000000", -- X := A, uPC := 0
   -- TXA
   b"0001_1000_0000_0_00_00_0011_00000000", -- A := X, uPC := 0
   -- TAY
   b"0000_0111_1001_0_00_00_0011_00000000", -- Y := A, uPC := 0
   -- TYA
   b"0001_1001_0000_0_00_00_0000_00000000", -- A := Y, uPC := 0
   -- ADC
   b"0100_0010_0000_0_00_00_0011_00000000", -- A += PM, uPC := 0
   -- SBC
   b"0101_0010_0000_0_00_00_0011_00000000", -- A -= PM, uPC := 0
   -- AND
   b"0110_0010_0000_0_00_00_0011_00000000", -- A := A AND PM, uPC := 0
   -- ORA
   b"0111_0010_0000_0_00_00_0011_00000000", -- A := A OR PM, uPC := 0
   -- EOR
   b"1000_0010_0000_0_00_00_0011_00000000", -- A := A XOR PM, uPC := 0
   -- ASL
   b"0000_0010_0000_0_10_00_0000_00000000", -- LC := PM
   b"0000_0000_0000_0_00_00_1100_00000000", -- uPC := 0 if LC = 0
   b"1010_0000_0000_0_01_00_1111_00000000", -- A := A << 1, LC--, uPC--
   -- LSR
   b"0000_0010_0000_0_10_00_0000_00000000", -- LC := PM
   b"0000_0000_0000_0_00_00_1100_00000000", -- uPC := 0 if LC = 0
   b"1100_0000_0000_0_01_00_1111_00000000", -- A := A << 1, LC--, uPC--
   -- INX
   b"0000_1010_1000_0_00_00_0011_00000000", -- X := X + 1, uPC := 0
   -- DEX
   b"0000_1011_1000_0_00_00_0011_00000000", -- X := X - 1, uPC := 0
   -- JMP
   b"0000_0010_0011_0_00_00_0011_00000000", -- PC := PM, uPC := 0
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000"
   );

signal u_mem : u_mem_t := u_mem_c;

begin  -- Behavioral
  uData <= u_mem(to_integer(uAddr));

end Behavioral;
