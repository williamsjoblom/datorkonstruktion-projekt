library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

-- pMem interface
entity pMem is
  port(
    pAddr : in unsigned(14 downto 0);
    pData : out unsigned(15 downto 0));
end pMem;

architecture Behavioral of pMem is

-- program Memory
type p_mem_t is array (0 to 4095) of unsigned(7 downto 0);
constant p_mem_c : p_mem_t := 
(
 x"9d"
,x"68"
,x"e0"
,x"9d"
,x"0f"
,x"e0"
,x"9d"
,x"d7"
,x"e3"
,x"9d"
,x"1e"
,x"e7"
,x"7d"
,x"09"
,x"e0"
,x"9d"
,x"55"
,x"e0"
,x"e0"
,x"06"
,x"e8"
,x"00"
,x"9d"
,x"22"
,x"e0"
,x"e0"
,x"0d"
,x"e8"
,x"0c"
,x"9d"
,x"22"
,x"e0"
,x"a0"
,x"00"
,x"9d"
,x"5e"
,x"e0"
,x"f1"
,x"13"
,x"20"
,x"9d"
,x"5e"
,x"e0"
,x"f9"
,x"13"
,x"20"
,x"a0"
,x"00"
,x"e0"
,x"08"
,x"9d"
,x"22"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"09"
,x"9d"
,x"22"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"0a"
,x"9d"
,x"22"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"07"
,x"9d"
,x"22"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"07"
,x"e8"
,x"f8"
,x"9d"
,x"22"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"07"
,x"e8"
,x"ff"
,x"9d"
,x"22"
,x"e0"
,x"a0"
,x"00"
,x"09"
,x"15"
,x"20"
,x"a8"
,x"01"
,x"cd"
,x"5e"
,x"e0"
,x"a0"
,x"00"
,x"08"
,x"00"
,x"81"
,x"02"
,x"20"
,x"81"
,x"03"
,x"20"
,x"a0"
,x"00"
,x"82"
,x"40"
,x"fa"
,x"41"
,x"18"
,x"00"
,x"20"
,x"00"
,x"e0"
,x"00"
,x"0f"
,x"40"
,x"00"
,x"a8"
,x"00"
,x"bd"
,x"8c"
,x"e0"
,x"9d"
,x"8e"
,x"e0"
,x"68"
,x"00"
,x"7d"
,x"7c"
,x"e0"
,x"a0"
,x"00"
,x"84"
,x"04"
,x"20"
,x"fc"
,x"06"
,x"20"
,x"9d"
,x"be"
,x"e0"
,x"a0"
,x"00"
,x"88"
,x"00"
,x"60"
,x"04"
,x"9d"
,x"a9"
,x"e0"
,x"90"
,x"00"
,x"40"
,x"0f"
,x"9d"
,x"a9"
,x"e0"
,x"a0"
,x"00"
,x"e8"
,x"f0"
,x"a8"
,x"0a"
,x"d5"
,x"b7"
,x"e0"
,x"30"
,x"30"
,x"9d"
,x"8e"
,x"e0"
,x"a0"
,x"00"
,x"30"
,x"37"
,x"9d"
,x"8e"
,x"e0"
,x"a0"
,x"00"
,x"09"
,x"02"
,x"20"
,x"a8"
,x"4f"
,x"bd"
,x"cd"
,x"e0"
,x"30"
,x"01"
,x"81"
,x"02"
,x"20"
,x"a0"
,x"00"
,x"08"
,x"00"
,x"81"
,x"02"
,x"20"
,x"09"
,x"03"
,x"20"
,x"a8"
,x"3b"
,x"bd"
,x"e1"
,x"e0"
,x"30"
,x"01"
,x"81"
,x"03"
,x"20"
,x"a0"
,x"00"
,x"08"
,x"00"
,x"81"
,x"03"
,x"20"
,x"a0"
,x"00"
,x"f1"
,x"02"
,x"20"
,x"f9"
,x"03"
,x"20"
,x"a0"
,x"00"
,x"43"
,x"68"
,x"20"
,x"41"
,x"20"
,x"20"
,x"20"
,x"20"
,x"43"
,x"68"
,x"20"
,x"42"
,x"20"
,x"20"
,x"20"
,x"20"
,x"43"
,x"68"
,x"20"
,x"43"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"00"
,x"20"
,x"28"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"29"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"29"
,x"20"
,x"20"
,x"28"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"29"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"29"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"2a"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"00"
,x"20"
,x"29"
,x"5c"
,x"20"
,x"29"
,x"20"
,x"20"
,x"28"
,x"20"
,x"2f"
,x"28"
,x"20"
,x"20"
,x"20"
,x"28"
,x"20"
,x"2f"
,x"28"
,x"20"
,x"20"
,x"29"
,x"5c"
,x"20"
,x"29"
,x"20"
,x"20"
,x"20"
,x"28"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"20"
,x"28"
,x"20"
,x"20"
,x"20"
,x"28"
,x"20"
,x"2f"
,x"28"
,x"20"
,x"20"
,x"20"
,x"28"
,x"20"
,x"2f"
,x"28"
,x"20"
,x"20"
,x"20"
,x"28"
,x"20"
,x"20"
,x"60"
,x"20"
,x"20"
,x"20"
,x"20"
,x"00"
,x"28"
,x"28"
,x"29"
,x"2f"
,x"28"
,x"20"
,x"20"
,x"29"
,x"5c"
,x"28"
,x"29"
,x"29"
,x"20"
,x"20"
,x"29"
,x"5c"
,x"28"
,x"29"
,x"29"
,x"28"
,x"28"
,x"29"
,x"2f"
,x"28"
,x"20"
,x"20"
,x"20"
,x"29"
,x"5c"
,x"20"
,x"20"
,x"20"
,x"20"
,x"28"
,x"20"
,x"29"
,x"5c"
,x"20"
,x"20"
,x"29"
,x"5c"
,x"28"
,x"29"
,x"29"
,x"20"
,x"20"
,x"29"
,x"5c"
,x"28"
,x"29"
,x"29"
,x"20"
,x"20"
,x"29"
,x"5c"
,x"29"
,x"29"
,x"28"
,x"20"
,x"20"
,x"20"
,x"00"
,x"20"
,x"2f"
,x"28"
,x"5f"
,x"29"
,x"29"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"5c"
,x"20"
,x"20"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"5c"
,x"20"
,x"20"
,x"2f"
,x"28"
,x"5f"
,x"29"
,x"29"
,x"28"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"20"
,x"20"
,x"20"
,x"29"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"5c"
,x"20"
,x"20"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"5c"
,x"20"
,x"20"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"28"
,x"29"
,x"5c"
,x"20"
,x"20"
,x"00"
,x"28"
,x"5f"
,x"29"
,x"29"
,x"20"
,x"20"
,x"20"
,x"20"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"20"
,x"20"
,x"5f"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"28"
,x"5f"
,x"29"
,x"29"
,x"20"
,x"20"
,x"29"
,x"5c"
,x"5f"
,x"5f"
,x"5f"
,x"20"
,x"20"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"5f"
,x"20"
,x"20"
,x"20"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"20"
,x"20"
,x"20"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"20"
,x"28"
,x"5f"
,x"28"
,x"29"
,x"28"
,x"28"
,x"5f"
,x"29"
,x"20"
,x"00"
,x"2f"
,x"20"
,x"5f"
,x"5f"
,x"7c"
,x"20"
,x"20"
,x"2f"
,x"20"
,x"5f"
,x"20"
,x"5c"
,x"20"
,x"7c"
,x"20"
,x"5c"
,x"7c"
,x"20"
,x"7c"
,x"7c"
,x"5f"
,x"20"
,x"5f"
,x"7c"
,x"28"
,x"28"
,x"2f"
,x"20"
,x"5f"
,x"5f"
,x"7c"
,x"20"
,x"20"
,x"7c"
,x"20"
,x"5f"
,x"20"
,x"29"
,x"20"
,x"2f"
,x"20"
,x"5f"
,x"20"
,x"5c"
,x"20"
,x"20"
,x"2f"
,x"20"
,x"5f"
,x"20"
,x"5c"
,x"20"
,x"7c"
,x"20"
,x"20"
,x"5c"
,x"2f"
,x"20"
,x"20"
,x"7c"
,x"20"
,x"00"
,x"5c"
,x"5f"
,x"5f"
,x"20"
,x"5c"
,x"20"
,x"7c"
,x"20"
,x"28"
,x"5f"
,x"29"
,x"20"
,x"7c"
,x"7c"
,x"20"
,x"2e"
,x"60"
,x"20"
,x"7c"
,x"20"
,x"7c"
,x"20"
,x"7c"
,x"20"
,x"20"
,x"7c"
,x"20"
,x"28"
,x"5f"
,x"5f"
,x"20"
,x"20"
,x"20"
,x"7c"
,x"20"
,x"5f"
,x"20"
,x"5c"
,x"7c"
,x"20"
,x"28"
,x"5f"
,x"29"
,x"20"
,x"7c"
,x"7c"
,x"20"
,x"28"
,x"5f"
,x"29"
,x"20"
,x"7c"
,x"7c"
,x"20"
,x"7c"
,x"5c"
,x"2f"
,x"7c"
,x"20"
,x"7c"
,x"20"
,x"00"
,x"7c"
,x"5f"
,x"5f"
,x"5f"
,x"2f"
,x"20"
,x"20"
,x"5c"
,x"5f"
,x"5f"
,x"5f"
,x"2f"
,x"20"
,x"7c"
,x"5f"
,x"7c"
,x"5c"
,x"5f"
,x"7c"
,x"7c"
,x"5f"
,x"5f"
,x"5f"
,x"7c"
,x"20"
,x"20"
,x"5c"
,x"5f"
,x"5f"
,x"5f"
,x"7c"
,x"20"
,x"20"
,x"7c"
,x"5f"
,x"5f"
,x"5f"
,x"2f"
,x"20"
,x"5c"
,x"5f"
,x"5f"
,x"5f"
,x"2f"
,x"20"
,x"20"
,x"5c"
,x"5f"
,x"5f"
,x"5f"
,x"2f"
,x"20"
,x"7c"
,x"5f"
,x"7c"
,x"20"
,x"20"
,x"7c"
,x"5f"
,x"7c"
,x"20"
,x"00"
,x"4b"
,x"65"
,x"79"
,x"20"
,x"3a"
,x"20"
,x"4e"
,x"6f"
,x"74"
,x"65"
,x"00"
,x"20"
,x"20"
,x"31"
,x"20"
,x"3a"
,x"20"
,x"43"
,x"00"
,x"20"
,x"20"
,x"32"
,x"20"
,x"3a"
,x"20"
,x"43"
,x"23"
,x"00"
,x"20"
,x"20"
,x"33"
,x"20"
,x"3a"
,x"20"
,x"44"
,x"00"
,x"20"
,x"20"
,x"34"
,x"20"
,x"3a"
,x"20"
,x"44"
,x"23"
,x"00"
,x"20"
,x"20"
,x"35"
,x"20"
,x"3a"
,x"20"
,x"45"
,x"00"
,x"20"
,x"20"
,x"36"
,x"20"
,x"3a"
,x"20"
,x"46"
,x"00"
,x"20"
,x"20"
,x"37"
,x"20"
,x"3a"
,x"20"
,x"46"
,x"23"
,x"00"
,x"20"
,x"20"
,x"38"
,x"20"
,x"3a"
,x"20"
,x"47"
,x"00"
,x"20"
,x"20"
,x"39"
,x"20"
,x"3a"
,x"20"
,x"47"
,x"23"
,x"00"
,x"20"
,x"20"
,x"41"
,x"20"
,x"3a"
,x"20"
,x"41"
,x"00"
,x"20"
,x"20"
,x"42"
,x"20"
,x"3a"
,x"20"
,x"41"
,x"23"
,x"00"
,x"20"
,x"20"
,x"43"
,x"20"
,x"3a"
,x"20"
,x"42"
,x"00"
,x"20"
,x"46"
,x"46"
,x"20"
,x"3a"
,x"20"
,x"6d"
,x"75"
,x"74"
,x"65"
,x"00"
,x"43"
,x"20"
,x"00"
,x"43"
,x"23"
,x"00"
,x"44"
,x"20"
,x"00"
,x"44"
,x"23"
,x"00"
,x"45"
,x"20"
,x"00"
,x"46"
,x"20"
,x"00"
,x"46"
,x"23"
,x"00"
,x"47"
,x"20"
,x"00"
,x"47"
,x"23"
,x"00"
,x"41"
,x"20"
,x"00"
,x"41"
,x"23"
,x"00"
,x"42"
,x"20"
,x"00"
,x"2d"
,x"2d"
,x"20"
,x"00"
,x"65"
,x"72"
,x"00"
,x"08"
,x"00"
,x"82"
,x"60"
,x"82"
,x"61"
,x"08"
,x"01"
,x"82"
,x"6d"
,x"e8"
,x"0f"
,x"9d"
,x"30"
,x"e0"
,x"9d"
,x"37"
,x"e0"
,x"9d"
,x"3e"
,x"e0"
,x"9d"
,x"70"
,x"e8"
,x"e0"
,x"0b"
,x"e8"
,x"e0"
,x"08"
,x"f0"
,x"9d"
,x"72"
,x"e0"
,x"9d"
,x"f9"
,x"e7"
,x"9d"
,x"11"
,x"e8"
,x"9d"
,x"29"
,x"e8"
,x"e0"
,x"00"
,x"e8"
,x"01"
,x"9d"
,x"e8"
,x"e0"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"9d"
,x"f4"
,x"e4"
,x"a0"
,x"00"
,x"e0"
,x"14"
,x"e8"
,x"01"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"f0"
,x"e8"
,x"e3"
,x"08"
,x"31"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"14"
,x"e8"
,x"02"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"f0"
,x"e8"
,x"e3"
,x"08"
,x"3c"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"14"
,x"e8"
,x"03"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"f0"
,x"e8"
,x"e3"
,x"08"
,x"44"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"14"
,x"e8"
,x"04"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"f0"
,x"e8"
,x"e3"
,x"08"
,x"4d"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"14"
,x"e8"
,x"05"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"f0"
,x"e8"
,x"e3"
,x"08"
,x"55"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"14"
,x"e8"
,x"06"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"f0"
,x"e8"
,x"e3"
,x"08"
,x"5e"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"14"
,x"e8"
,x"07"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"f0"
,x"e8"
,x"e3"
,x"08"
,x"66"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"14"
,x"e8"
,x"08"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"f0"
,x"e8"
,x"e3"
,x"08"
,x"6e"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"14"
,x"e8"
,x"09"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"f0"
,x"e8"
,x"e3"
,x"08"
,x"77"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"14"
,x"e8"
,x"0a"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"f0"
,x"e8"
,x"e3"
,x"08"
,x"7f"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"14"
,x"e8"
,x"0b"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"f0"
,x"e8"
,x"e3"
,x"08"
,x"88"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"14"
,x"e8"
,x"0c"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"f0"
,x"e8"
,x"e3"
,x"08"
,x"90"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"14"
,x"e8"
,x"0d"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"f0"
,x"e8"
,x"e3"
,x"08"
,x"99"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"14"
,x"e8"
,x"0e"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"f0"
,x"e8"
,x"e3"
,x"08"
,x"a1"
,x"9d"
,x"72"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"09"
,x"e8"
,x"29"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"e0"
,x"e8"
,x"e1"
,x"08"
,x"41"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"09"
,x"e8"
,x"2a"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"e0"
,x"e8"
,x"e1"
,x"08"
,x"7f"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"09"
,x"e8"
,x"2b"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"e0"
,x"e8"
,x"e1"
,x"08"
,x"bd"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"09"
,x"e8"
,x"2c"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"e0"
,x"e8"
,x"e1"
,x"08"
,x"fb"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"09"
,x"e8"
,x"2d"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"e0"
,x"e8"
,x"e2"
,x"08"
,x"39"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"09"
,x"e8"
,x"2e"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"f0"
,x"e8"
,x"e2"
,x"08"
,x"77"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"09"
,x"e8"
,x"2f"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"f0"
,x"e8"
,x"e2"
,x"08"
,x"b5"
,x"9d"
,x"72"
,x"e0"
,x"e0"
,x"09"
,x"e8"
,x"30"
,x"9d"
,x"e8"
,x"e0"
,x"e0"
,x"f0"
,x"e8"
,x"e2"
,x"08"
,x"f3"
,x"9d"
,x"72"
,x"e0"
,x"a0"
,x"00"
,x"e8"
,x"f8"
,x"fa"
,x"6c"
,x"9d"
,x"45"
,x"e0"
,x"a0"
,x"00"
,x"e8"
,x"ff"
,x"fa"
,x"6c"
,x"9d"
,x"45"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"6c"
,x"40"
,x"fe"
,x"82"
,x"6c"
,x"20"
,x"00"
,x"9d"
,x"45"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"6c"
,x"40"
,x"fd"
,x"82"
,x"6c"
,x"20"
,x"00"
,x"9d"
,x"45"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"6c"
,x"40"
,x"fb"
,x"82"
,x"6c"
,x"20"
,x"00"
,x"9d"
,x"45"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"6c"
,x"48"
,x"01"
,x"82"
,x"6c"
,x"20"
,x"00"
,x"9d"
,x"45"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"6c"
,x"48"
,x"02"
,x"82"
,x"6c"
,x"20"
,x"00"
,x"9d"
,x"45"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"6c"
,x"48"
,x"04"
,x"82"
,x"6c"
,x"20"
,x"00"
,x"9d"
,x"45"
,x"e0"
,x"a0"
,x"00"
,x"09"
,x"08"
,x"20"
,x"40"
,x"08"
,x"a8"
,x"00"
,x"bd"
,x"ed"
,x"e5"
,x"09"
,x"08"
,x"20"
,x"40"
,x"08"
,x"a8"
,x"00"
,x"cd"
,x"e0"
,x"e5"
,x"9d"
,x"78"
,x"e6"
,x"09"
,x"08"
,x"20"
,x"40"
,x"04"
,x"a8"
,x"00"
,x"bd"
,x"04"
,x"e6"
,x"09"
,x"08"
,x"20"
,x"40"
,x"04"
,x"a8"
,x"00"
,x"cd"
,x"f7"
,x"e5"
,x"9d"
,x"8d"
,x"e6"
,x"09"
,x"08"
,x"20"
,x"40"
,x"02"
,x"a8"
,x"00"
,x"bd"
,x"1b"
,x"e6"
,x"09"
,x"08"
,x"20"
,x"40"
,x"02"
,x"a8"
,x"00"
,x"cd"
,x"0e"
,x"e6"
,x"9d"
,x"a2"
,x"e6"
,x"09"
,x"08"
,x"20"
,x"40"
,x"01"
,x"a8"
,x"00"
,x"bd"
,x"32"
,x"e6"
,x"09"
,x"08"
,x"20"
,x"40"
,x"01"
,x"a8"
,x"00"
,x"cd"
,x"25"
,x"e6"
,x"9d"
,x"b7"
,x"e6"
,x"a0"
,x"00"
,x"9d"
,x"48"
,x"e6"
,x"0a"
,x"60"
,x"58"
,x"03"
,x"10"
,x"00"
,x"0a"
,x"61"
,x"30"
,x"01"
,x"20"
,x"00"
,x"9d"
,x"e8"
,x"e0"
,x"a0"
,x"00"
,x"0a"
,x"61"
,x"a8"
,x"00"
,x"d5"
,x"56"
,x"e6"
,x"08"
,x"26"
,x"82"
,x"61"
,x"7d"
,x"5f"
,x"e6"
,x"a8"
,x"27"
,x"c5"
,x"5f"
,x"e6"
,x"08"
,x"00"
,x"82"
,x"61"
,x"0a"
,x"60"
,x"a8"
,x"00"
,x"d5"
,x"6d"
,x"e6"
,x"08"
,x"02"
,x"82"
,x"60"
,x"7d"
,x"76"
,x"e6"
,x"a8"
,x"03"
,x"c5"
,x"76"
,x"e6"
,x"08"
,x"00"
,x"82"
,x"60"
,x"a0"
,x"00"
,x"08"
,x"f0"
,x"84"
,x"06"
,x"20"
,x"0a"
,x"61"
,x"38"
,x"01"
,x"82"
,x"61"
,x"9d"
,x"34"
,x"e6"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"08"
,x"f0"
,x"84"
,x"06"
,x"20"
,x"0a"
,x"60"
,x"30"
,x"01"
,x"82"
,x"60"
,x"9d"
,x"34"
,x"e6"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"08"
,x"f0"
,x"84"
,x"06"
,x"20"
,x"0a"
,x"61"
,x"30"
,x"01"
,x"82"
,x"61"
,x"9d"
,x"34"
,x"e6"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"9d"
,x"88"
,x"e8"
,x"a0"
,x"00"
,x"08"
,x"f0"
,x"84"
,x"06"
,x"20"
,x"0a"
,x"60"
,x"38"
,x"01"
,x"82"
,x"60"
,x"9d"
,x"34"
,x"e6"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"9d"
,x"6a"
,x"e9"
,x"a8"
,x"01"
,x"bd"
,x"db"
,x"e6"
,x"a0"
,x"00"
,x"9d"
,x"4f"
,x"e9"
,x"a8"
,x"01"
,x"c5"
,x"db"
,x"e6"
,x"58"
,x"04"
,x"82"
,x"6f"
,x"9d"
,x"4f"
,x"e9"
,x"4a"
,x"6f"
,x"20"
,x"00"
,x"e2"
,x"61"
,x"0a"
,x"60"
,x"a8"
,x"00"
,x"bd"
,x"01"
,x"e7"
,x"a8"
,x"01"
,x"bd"
,x"0a"
,x"e7"
,x"a8"
,x"02"
,x"bd"
,x"13"
,x"e7"
,x"fb"
,x"00"
,x"10"
,x"9d"
,x"f9"
,x"e7"
,x"7d"
,x"19"
,x"e7"
,x"fb"
,x"00"
,x"11"
,x"9d"
,x"11"
,x"e8"
,x"7d"
,x"19"
,x"e7"
,x"fb"
,x"00"
,x"12"
,x"9d"
,x"29"
,x"e8"
,x"9d"
,x"34"
,x"e6"
,x"a0"
,x"00"
,x"9d"
,x"d6"
,x"e5"
,x"9d"
,x"d1"
,x"e6"
,x"a0"
,x"00"
,x"a8"
,x"ff"
,x"bd"
,x"3d"
,x"e7"
,x"88"
,x"00"
,x"60"
,x"04"
,x"9d"
,x"a9"
,x"e0"
,x"90"
,x"00"
,x"e0"
,x"f0"
,x"40"
,x"0f"
,x"9d"
,x"48"
,x"e7"
,x"a0"
,x"00"
,x"e0"
,x"f0"
,x"e8"
,x"e3"
,x"08"
,x"d0"
,x"9d"
,x"72"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"00"
,x"cd"
,x"56"
,x"e7"
,x"e8"
,x"e3"
,x"08"
,x"ac"
,x"9d"
,x"72"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"01"
,x"cd"
,x"64"
,x"e7"
,x"e8"
,x"e3"
,x"08"
,x"af"
,x"9d"
,x"72"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"02"
,x"cd"
,x"72"
,x"e7"
,x"e8"
,x"e3"
,x"08"
,x"b2"
,x"9d"
,x"72"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"03"
,x"cd"
,x"80"
,x"e7"
,x"e8"
,x"e3"
,x"08"
,x"b5"
,x"9d"
,x"72"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"04"
,x"cd"
,x"8e"
,x"e7"
,x"e8"
,x"e3"
,x"08"
,x"b8"
,x"9d"
,x"72"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"05"
,x"cd"
,x"9c"
,x"e7"
,x"e8"
,x"e3"
,x"08"
,x"bb"
,x"9d"
,x"72"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"06"
,x"cd"
,x"aa"
,x"e7"
,x"e8"
,x"e3"
,x"08"
,x"be"
,x"9d"
,x"72"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"07"
,x"cd"
,x"b8"
,x"e7"
,x"e8"
,x"e3"
,x"08"
,x"c1"
,x"9d"
,x"72"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"08"
,x"cd"
,x"c6"
,x"e7"
,x"e8"
,x"e3"
,x"08"
,x"c4"
,x"9d"
,x"72"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"09"
,x"cd"
,x"d4"
,x"e7"
,x"e8"
,x"e3"
,x"08"
,x"c7"
,x"9d"
,x"72"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"0a"
,x"cd"
,x"e2"
,x"e7"
,x"e8"
,x"e3"
,x"08"
,x"ca"
,x"9d"
,x"72"
,x"e0"
,x"a0"
,x"00"
,x"a8"
,x"0b"
,x"cd"
,x"f0"
,x"e7"
,x"e8"
,x"e3"
,x"08"
,x"cd"
,x"9d"
,x"72"
,x"e0"
,x"a0"
,x"00"
,x"e8"
,x"e3"
,x"08"
,x"d4"
,x"9d"
,x"72"
,x"e0"
,x"a0"
,x"00"
,x"e0"
,x"00"
,x"e8"
,x"01"
,x"9d"
,x"e8"
,x"e0"
,x"e8"
,x"10"
,x"08"
,x"00"
,x"9d"
,x"41"
,x"e8"
,x"9d"
,x"34"
,x"e6"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"e0"
,x"08"
,x"e8"
,x"01"
,x"9d"
,x"e8"
,x"e0"
,x"e8"
,x"11"
,x"08"
,x"00"
,x"9d"
,x"41"
,x"e8"
,x"9d"
,x"34"
,x"e6"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"e0"
,x"10"
,x"e8"
,x"01"
,x"9d"
,x"e8"
,x"e0"
,x"e8"
,x"12"
,x"08"
,x"00"
,x"9d"
,x"41"
,x"e8"
,x"9d"
,x"34"
,x"e6"
,x"08"
,x"0f"
,x"84"
,x"06"
,x"20"
,x"a0"
,x"00"
,x"82"
,x"50"
,x"fa"
,x"51"
,x"e0"
,x"00"
,x"18"
,x"00"
,x"88"
,x"00"
,x"0f"
,x"50"
,x"00"
,x"9d"
,x"26"
,x"e7"
,x"90"
,x"00"
,x"10"
,x"00"
,x"09"
,x"02"
,x"20"
,x"38"
,x"03"
,x"81"
,x"02"
,x"20"
,x"09"
,x"03"
,x"20"
,x"30"
,x"01"
,x"81"
,x"03"
,x"20"
,x"68"
,x"00"
,x"18"
,x"00"
,x"a8"
,x"27"
,x"cd"
,x"47"
,x"e8"
,x"a0"
,x"00"
,x"e0"
,x"00"
,x"08"
,x"ff"
,x"83"
,x"00"
,x"10"
,x"83"
,x"00"
,x"11"
,x"83"
,x"00"
,x"12"
,x"68"
,x"00"
,x"18"
,x"00"
,x"a8"
,x"27"
,x"cd"
,x"72"
,x"e8"
,x"a0"
,x"00"
,x"08"
,x"00"
,x"88"
,x"00"
,x"9d"
,x"76"
,x"e5"
,x"90"
,x"00"
,x"10"
,x"00"
,x"9d"
,x"08"
,x"e9"
,x"88"
,x"00"
,x"9d"
,x"c3"
,x"e8"
,x"90"
,x"00"
,x"10"
,x"00"
,x"88"
,x"00"
,x"9d"
,x"da"
,x"e8"
,x"90"
,x"00"
,x"10"
,x"00"
,x"88"
,x"00"
,x"9d"
,x"f1"
,x"e8"
,x"90"
,x"00"
,x"30"
,x"01"
,x"a8"
,x"27"
,x"bd"
,x"be"
,x"e8"
,x"88"
,x"00"
,x"9d"
,x"3b"
,x"e9"
,x"7d"
,x"8c"
,x"e8"
,x"9d"
,x"7f"
,x"e5"
,x"a0"
,x"00"
,x"e3"
,x"00"
,x"10"
,x"18"
,x"00"
,x"a8"
,x"ff"
,x"cd"
,x"d2"
,x"e8"
,x"9d"
,x"af"
,x"e5"
,x"a0"
,x"00"
,x"9d"
,x"5e"
,x"e0"
,x"f1"
,x"10"
,x"20"
,x"a0"
,x"00"
,x"e3"
,x"00"
,x"11"
,x"18"
,x"00"
,x"a8"
,x"ff"
,x"cd"
,x"e9"
,x"e8"
,x"9d"
,x"bc"
,x"e5"
,x"a0"
,x"00"
,x"9d"
,x"5e"
,x"e0"
,x"f1"
,x"11"
,x"20"
,x"a0"
,x"00"
,x"e3"
,x"00"
,x"12"
,x"18"
,x"00"
,x"a8"
,x"ff"
,x"cd"
,x"00"
,x"e9"
,x"9d"
,x"c9"
,x"e5"
,x"a0"
,x"00"
,x"9d"
,x"5e"
,x"e0"
,x"f1"
,x"12"
,x"20"
,x"a0"
,x"00"
,x"18"
,x"00"
,x"88"
,x"00"
,x"9d"
,x"30"
,x"e9"
,x"e8"
,x"f0"
,x"08"
,x"20"
,x"9d"
,x"8e"
,x"e0"
,x"90"
,x"00"
,x"88"
,x"00"
,x"10"
,x"00"
,x"30"
,x"01"
,x"82"
,x"6d"
,x"9d"
,x"30"
,x"e9"
,x"e8"
,x"f0"
,x"08"
,x"3c"
,x"9d"
,x"8e"
,x"e0"
,x"90"
,x"00"
,x"10"
,x"00"
,x"a0"
,x"00"
,x"0a"
,x"6d"
,x"20"
,x"00"
,x"e0"
,x"14"
,x"9d"
,x"e8"
,x"e0"
,x"a0"
,x"00"
,x"08"
,x"0a"
,x"e0"
,x"fa"
,x"88"
,x"00"
,x"9d"
,x"7c"
,x"e9"
,x"90"
,x"00"
,x"38"
,x"01"
,x"a8"
,x"00"
,x"cd"
,x"3f"
,x"e9"
,x"a0"
,x"00"
,x"09"
,x"09"
,x"20"
,x"40"
,x"f0"
,x"a8"
,x"00"
,x"cd"
,x"4f"
,x"e9"
,x"e1"
,x"09"
,x"20"
,x"09"
,x"09"
,x"20"
,x"40"
,x"f0"
,x"a8"
,x"00"
,x"bd"
,x"5c"
,x"e9"
,x"18"
,x"00"
,x"a0"
,x"00"
,x"09"
,x"09"
,x"20"
,x"40"
,x"f0"
,x"a8"
,x"00"
,x"bd"
,x"78"
,x"e9"
,x"08"
,x"00"
,x"a0"
,x"00"
,x"08"
,x"01"
,x"a0"
,x"00"
,x"e8"
,x"ff"
,x"28"
,x"00"
,x"38"
,x"01"
,x"20"
,x"00"
,x"a8"
,x"00"
,x"cd"
,x"7e"
,x"e9"
,x"18"
,x"00"
,x"38"
,x"01"
,x"10"
,x"00"
,x"a8"
,x"00"
,x"cd"
,x"7c"
,x"e9"
,x"a0"
,x"00"
,x"77"
,x"0b"
,x"a6"
,x"47"
,x"ec"
,x"97"
,x"47"
,x"fb"
,x"b3"
,x"70"
,x"30"
,x"f4"
,x"00"
,x"00"
,x"00"
,x"00"
,x"bb"
,x"85"
,x"53"
,x"23"
,x"f6"
,x"cb"
,x"a3"
,x"7d"
,x"59"
,x"38"
,x"18"
,x"fa"
,x"00"
,x"00"
,x"00"
,x"00"
,x"dd"
,x"c2"
,x"a9"
,x"91"
,x"7b"
,x"65"
,x"51"
,x"3e"
,x"2c"
,x"1c"
,x"0c"
,x"fd"
,x"00"
,x"00"
,x"00"
,x"00"
,x"ee"
,x"e1"
,x"d4"
,x"c8"
,x"bd"
,x"b2"
,x"a8"
,x"9f"
,x"96"
,x"8e"
,x"86"
,x"7e"
,x"00"
,x"00"
,x"00"
,x"00"
,x"77"
,x"70"
,x"6a"
,x"64"
,x"5e"
,x"59"
,x"54"
,x"4f"
,x"4b"
,x"47"
,x"43"
,x"3f"
,x"00"
,x"00"
,x"00"
,x"00"
,x"3b"
,x"38"
,x"35"
,x"32"
,x"2f"
,x"2c"
,x"2a"
,x"27"
,x"25"
,x"23"
,x"21"
,x"1f"
,x"00"
,x"00"
,x"00"
,x"00"
,x"1d"
,x"1c"
,x"1a"
,x"19"
,x"17"
,x"16"
,x"15"
,x"13"
,x"12"
,x"11"
,x"10"
,x"0f"
,x"00"
,x"00"
,x"00"
,x"00"
,x"0e"
,x"0e"
,x"0d"
,x"0c"
,x"0b"
,x"0b"
,x"0a"
,x"09"
,x"09"
,x"08"
,x"08"
,x"07"
,x"00"
,x"00"
,x"00"
,x"00"
,x"07"
,x"07"
,x"06"
,x"06"
,x"05"
,x"05"
,x"05"
,x"04"
,x"04"
,x"04"
,x"04"
,x"03"
,x"00"
,x"00"
,x"00"
,x"00"
,x"07"
,x"07"
,x"06"
,x"06"
,x"05"
,x"05"
,x"05"
,x"04"
,x"04"
,x"04"
,x"04"
,x"03"
,x"00"
,x"00"
,x"00"
,x"00"
,x"03"
,x"03"
,x"03"
,x"03"
,x"02"
,x"02"
,x"02"
,x"02"
,x"02"
,x"02"
,x"02"
,x"01"
,x"00"
,x"00"
,x"00"
,x"00"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"01"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"e0"
);


  signal p_mem : p_mem_t := p_mem_c;


begin  -- pMem
  pData <= p_mem(to_integer(pAddr(11 downto 0) + 1)) & p_mem(to_integer(pAddr(11 downto 0)));

end Behavioral;

