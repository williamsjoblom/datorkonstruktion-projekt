library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

-- uMem interface
entity uMem is
  port (
    uAddr : in unsigned(7 downto 0);
    uData : out unsigned(28 downto 0));
end uMem;

architecture Behavioral of uMem is


-- micro Memory
type u_mem_t is array (0 to 255) of unsigned(28 downto 0);
constant u_mem_c : u_mem_t :=
  -- ALU__TB___FB__PC_LC_ST_SEQ__uAddr
   -- Fetch
  (b"0000_0011_1110_0_00_00_0000_00000000", -- ASR := PC
   b"0000_0000_0000_1_00_00_0000_00000000", -- PC++
   b"0000_0010_0001_0_00_00_0000_00000000", -- IR := PM
   -- E-A Calculation
   b"0000_0000_0000_0_00_00_0010_00000000", -- uPC := K2
   -- Immediate Addressing: LDA #10
   b"0000_0011_1110_1_00_00_0000_00000000", -- ASR := PC, PC++
   b"0000_0000_0000_0_00_00_0001_00000000", -- uPC := K1
   -- Absolute Addressing: LDA $FF77
   b"0000_0011_1110_1_00_00_0000_00000000", -- ASR := PC, PC++
   b"0000_0000_0000_1_00_00_0000_00000000", -- PC++
   b"0000_0010_1110_0_00_00_0000_00000000", -- ASR := PM
   b"0000_0000_0000_0_00_00_0001_00000000", -- uPC := K1
   -- ZP Absolute Addressing: JMP $33
   b"0000_0011_1110_1_00_00_0000_00000000", -- ASR := PC, PC++
   b"0000_0000_0000_0_00_00_0000_00000000", -- NOP (wait for RAM)
   b"0000_0010_1110_0_00_00_0000_00000000", -- ASR := PM,
   b"0000_0000_1111_0_00_00_0000_00000000", -- ASRmsb := 0
   b"0000_0000_0000_0_00_00_0001_00000000", -- uPC := K1
   -- Absolute X: STA $AA16, X
   b"0000_0011_1110_1_00_00_0000_00000000", -- ASR := PC, PC++
   b"0000_0000_0000_1_00_00_0000_00000000", -- PC++
   b"0000_0010_1101_0_00_00_0000_00000000", -- ASR := PM[X]
   b"0000_0000_0000_0_00_00_0001_00000000", -- uPC := K1
   -- Indirect: ($300)
   b"0000_0011_1110_1_00_00_0000_00000000", -- ASR := PC, PC++
   b"0000_0000_0000_1_00_00_0000_00000000", -- PC++
   b"0000_0010_1110_0_00_00_0000_00000000", -- ASR := PM
   b"0000_0000_0000_0_00_00_0000_00000000", -- NOP (wait for RAM)
   b"0000_0010_1110_0_00_00_0000_00000000", -- ASR := PM
   b"0000_0000_0000_0_00_00_0001_00000000", -- uPC := K1
   -- Absolute Jump: JMP $1234
   b"0000_0011_1110_1_00_00_0000_00000000", -- ASR := PC, PC++
   b"0000_0000_0000_1_00_00_0001_00000000", -- PC++, uPC := K1

   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   -- Indexed Indirect X: ($1337, X)
   b"0000_0011_1110_1_00_00_0000_00000000", -- ASR := PC, PC++
   b"0000_0000_0000_1_00_00_0000_00000000", -- PC++
   b"0000_0010_1101_0_00_00_0000_00000000", -- ASR := PM[X]
   b"0000_0000_0000_0_00_00_0000_00000000", -- NOP (wait for RAM)
   b"0000_0010_1110_0_00_00_0000_00000000", -- ASR := PM
   b"0000_0000_0000_0_00_00_0001_00000000", -- uPC := K1
   -- Indirect Indexed X: ($1337), X
   b"0000_0011_1110_1_00_00_0000_00000000", -- ASR := PC, PC++
   b"0000_0000_0000_1_00_00_0000_00000000", -- PC++
   b"0000_0010_1110_0_00_00_0000_00000000", -- ASR := PM
   b"0000_0000_0000_0_00_00_0000_00000000", -- NOP (wait for RAM)
   b"0000_0010_1101_0_00_00_0000_00000000", -- ASR := PM[X]
   b"0000_0000_0000_0_00_00_0001_00000000", -- uPC := K1
   
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   -- NOP
   b"0000_0000_0000_0_00_00_0011_00000000", -- uPC := 0
   -- LDA
   b"0001_0010_0000_0_00_00_0011_00000000", -- A := PM, uPC := 0
   -- TAX
   b"0000_0111_1000_0_00_00_0011_00000000", -- X := A, uPC := 0
   -- TXA
   b"0001_1000_0000_0_00_00_0011_00000000", -- A := X, uPC := 0
   -- TAY
   b"0000_0111_1001_0_00_00_0011_00000000", -- Y := A, uPC := 0
   -- TYA
   b"0001_1001_0000_0_00_00_0000_00000000", -- A := Y, uPC := 0
   -- ADC
   b"0100_0010_0000_0_00_00_0011_00000000", -- A += PM, uPC := 0
   -- SBC
   b"0101_0010_0000_0_00_00_0011_00000000", -- A -= PM, uPC := 0
   -- AND
   b"0110_0010_0000_0_00_00_0011_00000000", -- A := A AND PM, uPC := 0
   -- ORA
   b"0111_0010_0000_0_00_00_0011_00000000", -- A := A OR PM, uPC := 0
   -- EOR
   b"1000_0010_0000_0_00_00_0011_00000000", -- A := A XOR PM, uPC := 0
   -- ASL
   b"0000_0010_0000_0_10_00_0000_00000000", -- LC := PM
   b"0000_0000_0000_0_00_00_1100_00000000", -- uPC := 0 if LC = 0
   b"1010_0000_0000_0_01_00_1111_00000000", -- A := A << 1, LC--, uPC--
   -- LSR
   b"0000_0010_0000_0_10_00_0000_00000000", -- LC := PM
   b"0000_0000_0000_0_00_00_1100_00000000", -- uPC := 0 if LC = 0
   b"1100_0000_0000_0_01_00_1111_00000000", -- A := A << 1, LC--, uPC--
   -- INX
   b"0000_1010_1000_0_00_00_0011_00000000", -- X := X + 1, uPC := 0
   -- DEX
   b"0000_1011_1000_0_00_00_0011_00000000", -- X := X - 1, uPC := 0
   -- JMP
   b"0000_0010_0011_0_00_00_0011_00000000", -- PC := PM, uPC := 0
   -- STA
   b"0000_0111_0010_0_00_00_0011_00000000", -- PM := A, uPC := 0
   -- PHA
   b"0000_0111_1100_0_00_10_0011_00000000", -- (SP) := A, SP--, uPC := 0
   -- PLA
   b"0000_0000_0000_0_00_01_0000_00000000", -- SP++
   b"0001_1100_0000_0_00_00_0011_00000000", -- A := (SP), uPC := 0
   -- JSR : Candidate for optimization
   b"0000_0000_0000_0_00_00_0000_00000000", -- PC++ nope
   b"0000_0000_0000_0_00_00_0000_00000000", -- PC++ nope
   b"0000_0100_1100_0_00_10_0000_00000000", -- (SP) := PC, SP--
   b"0000_0000_0000_0_00_00_0000_00000000", -- NOP (wait for RAM)
   b"0000_0011_1100_0_00_10_0000_00000000", -- (SP) := PCmsb, SP--
   b"0000_0010_0011_0_00_00_0011_00000000", -- PC := PM, uPC := 0
   b"0000_0000_0000_0_00_00_0000_00000000",
   -- RTS
   b"0000_0000_0000_0_00_01_0000_00000000", -- SP++
   b"0000_0000_0000_0_00_00_0000_00000000", -- NOP (wait for ram)
   b"0000_1100_0011_0_00_01_0011_00000000", -- PC := (SP), SP++, uPC := 0
   -- CMP
   b"1111_0010_0000_0_00_00_0011_00000000", -- A cmp PM, uPC := 0
   -- BCS
   b"0000_0000_0000_0_00_00_1010_01000110", -- uPC := JMP if C = 1
   b"0000_0000_0000_0_00_00_0011_00000000", -- uPC := 0
   -- BEQ
   b"0000_0000_0000_0_00_00_1000_01000110", -- uPC := JMP if Z = 1
   b"0000_0000_0000_0_00_00_0011_00000000", -- uPC := 0
   -- BMI
   b"0000_0000_0000_0_00_00_1001_01000110", -- uPC := JMP if S = 1
   b"0000_0000_0000_0_00_00_0011_00000000", -- uPC := 0
   -- BNE
   b"0000_0000_0000_0_00_00_1000_00000000", -- uPC := 0 if Z = 1
   b"0000_0000_0000_0_00_00_0101_01000110", -- uPC := JMP
   -- BPL
   b"0000_0000_0000_0_00_00_1001_00000000", -- uPC := 0 if S = 1
   b"0000_0000_0000_0_00_00_0101_01000110", -- uPC := JMP
   -- BIT
   b"0011_0010_0000_0_00_00_0011_00000000", -- Z := 1 if A[PM] = 0, uPC := 0
   -- LDX
   b"0000_0010_1000_0_00_00_0011_00000000", -- X := PM, uPC := 0
   -- LDY
   b"0000_0010_1001_0_00_00_0011_00000000", -- Y := PM, uPC := 0
   -- STX
   b"0000_1000_0010_0_00_00_0011_00000000", -- PM := A, uPC := 0
   -- STY
   b"0000_1001_0010_0_00_00_0011_00000000", -- PM := Y, uPC := 0
   b"0000_0000_0000_0_00_00_0000_00000000",

   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000",
   b"0000_0000_0000_0_00_00_0000_00000000"
   );

signal u_mem : u_mem_t := u_mem_c;

begin  -- Behavioral
  uData <= u_mem(to_integer(uAddr));

end Behavioral;
