library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

-- pMem interface
entity pMem is
  port(
    pAddr : in unsigned(14 downto 0);
    pData : out unsigned(15 downto 0));
end pMem;

architecture Behavioral of pMem is

-- program Memory
type p_mem_t is array (0 to 255) of unsigned(7 downto 0);
constant p_mem_c : p_mem_t := 
(
 x"9d"
,x"48"
,x"e0"
,x"e0"
,x"00"
,x"e8"
,x"71"
,x"9d"
,x"69"
,x"e0"
,x"e0"
,x"01"
,x"e8"
,x"02"
,x"9d"
,x"69"
,x"e0"
,x"e8"
,x"f0"
,x"e0"
,x"13"
,x"9d"
,x"bb"
,x"e0"
,x"e0"
,x"0f"
,x"9d"
,x"bb"
,x"e0"
,x"e0"
,x"0e"
,x"9d"
,x"bb"
,x"e0"
,x"e0"
,x"09"
,x"9d"
,x"bb"
,x"e0"
,x"e0"
,x"03"
,x"9d"
,x"bb"
,x"e0"
,x"e0"
,x"00"
,x"9d"
,x"bb"
,x"e0"
,x"e0"
,x"02"
,x"9d"
,x"bb"
,x"e0"
,x"e0"
,x"0f"
,x"9d"
,x"bb"
,x"e0"
,x"e0"
,x"0f"
,x"9d"
,x"bb"
,x"e0"
,x"e0"
,x"0d"
,x"9d"
,x"bb"
,x"e0"
,x"7d"
,x"45"
,x"e0"
,x"9d"
,x"71"
,x"e0"
,x"e0"
,x"06"
,x"e8"
,x"00"
,x"9d"
,x"69"
,x"e0"
,x"e0"
,x"07"
,x"e8"
,x"f8"
,x"9d"
,x"69"
,x"e0"
,x"e0"
,x"08"
,x"e8"
,x"0f"
,x"9d"
,x"69"
,x"e0"
,x"e0"
,x"09"
,x"e8"
,x"0f"
,x"9d"
,x"69"
,x"e0"
,x"a0"
,x"00"
,x"9d"
,x"8e"
,x"e0"
,x"9d"
,x"7e"
,x"e0"
,x"a0"
,x"00"
,x"08"
,x"00"
,x"81"
,x"01"
,x"20"
,x"9d"
,x"a8"
,x"e0"
,x"9d"
,x"9e"
,x"e0"
,x"a0"
,x"00"
,x"f9"
,x"00"
,x"20"
,x"08"
,x"fe"
,x"81"
,x"01"
,x"20"
,x"9d"
,x"a8"
,x"e0"
,x"9d"
,x"9e"
,x"e0"
,x"a0"
,x"00"
,x"f1"
,x"00"
,x"20"
,x"08"
,x"ff"
,x"81"
,x"01"
,x"20"
,x"9d"
,x"a8"
,x"e0"
,x"9d"
,x"9e"
,x"e0"
,x"a0"
,x"00"
,x"08"
,x"04"
,x"81"
,x"01"
,x"20"
,x"9d"
,x"a8"
,x"e0"
,x"a0"
,x"00"
,x"08"
,x"28"
,x"38"
,x"01"
,x"cd"
,x"aa"
,x"e0"
,x"a0"
,x"00"
,x"08"
,x"00"
,x"81"
,x"02"
,x"20"
,x"81"
,x"03"
,x"20"
,x"a0"
,x"00"
,x"f4"
,x"04"
,x"20"
,x"fc"
,x"06"
,x"20"
,x"9d"
,x"c6"
,x"e0"
,x"a0"
,x"00"
,x"09"
,x"02"
,x"20"
,x"a8"
,x"4f"
,x"bd"
,x"d5"
,x"e0"
,x"30"
,x"01"
,x"81"
,x"02"
,x"20"
,x"a0"
,x"00"
,x"08"
,x"00"
,x"81"
,x"02"
,x"20"
,x"09"
,x"03"
,x"20"
,x"a8"
,x"3b"
,x"bd"
,x"e9"
,x"e0"
,x"30"
,x"01"
,x"81"
,x"03"
,x"20"
,x"a0"
,x"00"
,x"08"
,x"00"
,x"81"
,x"03"
,x"20"
,x"a0"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"00"
,x"e0"
);


  signal p_mem : p_mem_t := p_mem_c;


begin  -- pMem
  pData <= p_mem(to_integer(pAddr(7 downto 0) + 1)) & p_mem(to_integer(pAddr(7 downto 0)));

end Behavioral;

